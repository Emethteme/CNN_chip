//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2017 ICLAB Fall Course
//   MID			
//   Author     : YiWei Chen (andychen.ee01@g2.nctu.edu.tw)
//
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v1.0
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`ifdef RTL
    `timescale 1ns/10ps
    `include "CNN.v"  
    `define DELAY 0
`define CYCLE_TIME 10
    `define MODE 0
`endif
`ifdef GATE
    `timescale 1ns/1ps
    `define DELAY 0
    `include "CNN_SYN.v"
`define CYCLE_TIME 10
    `define MODE 1
`endif
`ifdef POSIM
    `timescale 1ns/1ps
`define DELAY 5
    `include "CHIP.v"
`define CYCLE_TIME 20
    `define MODE 2
`endif

module PATTERN(
    // Output signals
    clk,
    rst_n,
    in_valid_1,
    in_valid_2,
    in_data,
    // Input signals
    out_valid,
    number_2,
    number_4,
    number_6
);

`protected
IdKi5SQV5DT^<OkYNf@=[he9Ud5D75oo6]jB\ibdj><eQF0Am5e^DlP\6>REZD3J
D2fRH<FDB;\kAi8pQ\E[8ZHdYMX[D>D0N3e@DS?@LCR1ZOTPDdRMf3TWS??GAjbq
OGBVE?YW;XWdb5fU\JlNn9;M9EGKAO=83LM[mBedf^Cob9?R<hTo5enqbl\G^lpd
Kkoa1qDLPZZG3G[\]1FRQdiOMqc>j1NFB7YgYF1dE5KKP>q=I]=lZk6i2IK<8CVV
`Lm12N2BUXq[PZ<>_UdNjWi>X;:JUd6EkCgC0`qUWInRhPZRTPkBj[meF:13UUIM
eR<KIQ08M^jp0RD8cmHRBk3D>fl^iXeW]b<b:`V@_:R;AP9dB87HpdUg;YJqY^WK
KB[KC>h0GhGhdQT0DTQqmZS0^L@99G56jGmQEE4N3UqYeH3Qn9RNeNLU:j^:7OM>
lpD^dO9CbeiZB]?QB9?C[GWYJTEZK=pbbX\RWCkR6A7hcIkX7lY0Pq`n@FDhpb4c
[0=?iIYdoeZ^hXC6fN^_k1XDXS>GobXUlqeaOJDlQQ6GY1lg0UKeBC8Vj:TBZdN<
p5an;^BoIVM8T^9TY2;e:O;0Lo:=fS`ORaQ7cBH:86bT?UXJoAF1ASke_[:Yd>md
=C==6gcMQphD5jkGCH?jMo<aajP[U>4nd8`WWi:Ie2fSPaKC0qkhG@=[a?@VJaBK
OL]AcDFkm0@<q7FlRKoYc@Nf3<k2:Ia8d:L3V`B1M8W=BQR81DWYKYh2`i74q0?S
bfD=n]?S\bGN?ad<;<gqJKc6=l4nCTSnO2ihW<MgVMYbic\\glD^p78OAlA;;agk
OLDCk@:fH<O5m@<9SU7=;c2Fe>QqFLi71nHC?F\2]k]2:>hH\No9EJ@Qq:7OR8^A
D]8mTJ_SL]\mF=m16O;J_jHqc6JRKH[D6VdjA1F385kn>PcgBnY9]34Da5D8gN?[
Xo0Xlgc=h8kmLNVY5d=Cm@=@;V@kqD^ZGY=8m7i1H?UMH86hd^O^ffCX?l5f38Z0
`kh6el1NZnGh\PX=nZmMDJ0C@ZOkLHj18qAL4nUh48BeCa<]Af[M?DFh`e@l[[Z^
k]KGYY01[<G?8_7:^@Zo_Ia\a@JBXR1ZeA71q?d6LKc^Q=AooQhEj62o>nN66__:
2ig<P7SUVEEeHCfbbNWNW46Wk;=3Oek;9l8LdF]miCD`9PL\lp<2a=0??0F1NmMH
bocJLfcK@7q2N2;j0WZ4Rf2@LTJYc=`S\\Tp8fK<S@MA4?[gW6F[h@U^ONA]3<31
C>U`dX@Wd\d6M=DBE697j[q=_PRFT6iCee52[:AfCH58CIZ?mpm^f81j;SWk`mR:
:`>BH:;d[qa;?Q0lL1X6_42l4=:L_D]1pF7Z9aaDbkNLoF9^AcIEWX4Uok]2OYJ5
6eUnD`L>:o;_O^C^p_YMLM?23aYV4jiI`k\5SULGqoDMD_R=C16p@jNB2E8QJ>N3
D7]HODmBCJ_dqFjE8H1Y`W]cSW51ZkC[W503LB?Hh6k`8Y6N<c2Kl`ke:bQqj?9T
X`\@o97SoRMjQNC\O7bUhcVBOae=8XnhZY^G4345DZi7hSef96fBFILMbRGh<o:3
XE9YOmlk\<3qGT<11EbN3D=3dMc:7LU@k::=ql>2dBQ`O;6V=2d;2o;43G_GgoY\
^Whh_b^NapZB=?PNh;Y>0HL@KEGL[^D3<\a<@IkMIQqkPXe^Xqo7;\:7qA5?UeaT
A<=J>eCHXSg>WgOjM`o=Dl[ccpO3n1:?qS]\Sk@EDgj>cNDb:PB5KaZP3R2facAh
fMXL1l5Qfe?lD]Z=LDJa_h8ed1UG@iD0E_@k@pTMAX9?>b<aNZ?gEKDn?0`Y@Ymk
Vlh2omhJBBN]6X?OeA3RZFQ1bBof\1kPE;X7;_T^Qdp7G2[^hpPkbA;=p[<Fh4ai
2Cl<_3blj5a45Si\hn4WNbeN;UdW?J`7k8YPYgh3TNHQ\IR`QkX6k]CMF_nS[X>8
7q\PM9S]8Y5Ce9SBfWKoURmem:IOiWaTN_HXBN;Z3:2>O;1fH\nk0@Hlmbb\B5XJ
BTK_GI@e;Rimhp13@Gc1qOEL`0_IAULQY1DC^OLc?hED\VVZe:5hdfm`kdW0=pnB
ZSF_<kNKQoZI=X_H6oeIm<R;@]o5QQSN\N^d1RZDVQ@Q[eGS`RQ2bX5e[@7Kba]P
^fp=Da1J4LCJ>^BG>_jW7:Qk?Fa?CZKe5^`TKLM=g\]QK=>2Dm1KM<dLX?WCE^G8
YR;7^HIJd2;gFZ@mIa5Ro8FW5dSbopMLDR[o0kQ:JQ9mWP:MSmNa:31fek?Vi9M3
8BqZ^f_;kld`^5K@^`?@TOTClI^`m?Q^3dgmQNhYcXLQ;3`N`COoHGRW7?e4FTV@
E:HUZ:QSM8T1X1`lhJo^n0k_YG<hmp5YOKNn;Wf6]G\mgU37?5LgbmReiBWMaDXR
L3L[GFc4PPXoWC089GD[k[^L[eBG?PS04YWRMR0MNC@3GcB`]]^c=S@<pG5>F1ho
SpY=98bCfd00TgHIeiK2<V;L`YE`_2AC8a@1bLnGj6p_V3ESULEnenCK?o^kfRZF
79BDPM5@PN@8PjDO3;iEIO;\R1<=Ej0]>:?nUYMBG]Xc`q=D4j:K;oFe6CI]?k:l
8A?=Ef@CF]WEaLXgcWnFelVVGTEIBco>BA3C^HA?nW>D`ec\`EO9pYh4KceVRTaC
k5407UVCE6lgCN9LAagiT57CfO_imRUFFji[S`IVDJ;CZCiR?1SQ;YOV`C4<8W6j
b7a42?N_^0AUVNQ]pW7hF:kjI=B5cdk6eo0]\XmnkYSP;lVPbo]V8U;Hj1]3cDof
PE>dF]iJAh;4WJPoEWWg[o^aV^SiE<Bb>6jNLe0Ado`;qCEk?Hmf8m50:oCgkBjB
0_od68Fi;]li7>UC2X3`R?8[H[kLY8:TfoEm_lad309FNCoZXj7:FE_9_h=QEeh6
CV7?Ub4Vp2PHHQN^Iq[A5b^6_F@J8UHV`Dn7Ym[]CoAVXSoQQ]kX\ZWo7^pcW4MK
lOld:WmAUQd3V?19b=acdh<@_QFBNT3adgRJ:]dLZHh=kkIFd[nCeL5<]?^;VgfF
1pBP20K<6SY43KfSD0MI?kW>YaS[=4V]bP1\<ThQEE3:H;Y]HX@WZW0[k8;1d@e:
o8V3i]m2IQhQAMm]6=nea0O=M<NBdaN][pjX1^3FP12jOaBLac0aLdfc<L1Q4ie4
NSY_33@Z^`m3\i;FTjiD8MlJcaKI`<KOfFKDF\IW`5lbKn6:DPg4:_UF[VM_TB7O
Vq6X^m4YgI^<3kjD::;GjliOj9lHRL;nWe<io2ZPnD[XX5<Xn8]I^kV:il]Vg71H
KpQ?fC[:<>BR5FT=:kRBX<@EH12;gP^0_NaK0@XkU_n1abBH63E4?X5kVI_OXO^a
^4TP7kgV`i;::dCG3U^N[M^?<kD=ch\T9qKhh]=NN>q_CJ:=ZXplN[Q^YG\L9HbW
:b?N;i4hAk<q=<J\P^>Bl[^2o_==_XbU0KdSoX15E@mBbG9^JQ\jU9Vik9PAS[:?
5Qb16gOkD;Ck4>JHQTmSDM^LaaHQlhBSD1cCCndFEc3g?@26WoAEqD37OIne\i2p
DN3gEEMoR;M\@MHh?Fle02[Q\5\\qa7ZQIggi^?M]CSF43DCBJF1HDAg9PA^Nb2A
GQ::gpmJPfLa68RJEhN0XCFh6:;e[JoFaq<YNK7l<4LfjhT]O]aCU:[h`N0JM9pA
U0_ZU<]4Pa2QYM^BonQ\mpSf=<aIH`HgYYPlf\\=oQAOp3bA=G2EKq9W[2DHq0R8
l>3:0e3hlf@2@Th?HjnK[meZSh_h`Eo;T7==pW3:?N^YE0[RDJd[742X5c^QDTEh
Gh7hK6kOeENWq8]gX<SEnE_NRe1HeV^gkg^YbgU\JMBk>iE1O1^Jgc@Rb<Q^T[UN
bDQk;[GB95UXEqAi5]JQjXiBWNdf\0Vejo_NeckIVSJW6lBmS5m9@p_JNjX9QqYZ
HTV@nlE:iH:VAE9FRecg?08]YOhf\Sqnjg7kSApiWhRjL``FKI[=QV6H8hlqB`@G
36;pXhAODKpBioc\^RUne@ah8Gc`ef1ABjfKU>qK1WndJ6T@;Lg94[Q2@R\7;U?S
2N7jJUSaQY@ElqV\`ln0N[P1QX_DFJja`\93`8GNJIAA^0:N<qhA5HFb?qAe0FoL
=hlkBjZZ8b3ME@phL]8J8`@k\H]jP`F<5X1O7E1]SH0F\9GB^pHo9>IT12Lb9cQ0
gVNIPIp:_Pa?VBPBMg0HWA0JOiC:fMSHWRdoNi4f0]L<l:O4EXLkA0J1A2:>FlZ3
c?hc__5:KZ0naGDeIdm[T__ClFDnMHVYE[M1[9QQ364_mPL@8<ML_YC0Ip9MkV94
YHDK`kZdk4VO>LR:Mhm`m[>Wc6??Yja2dWO0G>El7f>VP0`3gWO_;:5^lLfBb_N:
On_lHfaF9bk;2b9TPq4DKll;L28PD7Wl[:?FD@XDH<R:BoNbPZSj^XN_3?nnDPFR
Bj?=7^X:Aj<kXJcGRo44Rkd6?_8cli`haA_9Dadn`qAl[MVIXT_a:Q9k_2<<m:4_
OV_gA]KV9\l9C@iR5\89inN>M:_T50VmATH1qOb_37A4g`\I<E8W_<NK9cPKl16l
oaTGCoLjVQA\0MXj2mIFhU=9No>Aim]BD8\EAIf3j@IDcTLRR9D5\dNN4M04^GYI
X?94i9oTDPUQbp0dIdLdTFDJeITda3hPeh?@cQG^3oM4JP9OU<<955H7N_H5lAdj
=neA;gdNe^=4dELm06<GQ<hBm_oWFoVE:]W;:qGQX302UoGgGY;?k331pWS10N]h
FOQ@cclpVN:SBHM;Y^H:^kTU49pbFdblcb<qI1W]\j`qUMlUXEO5ma=nmZMN@S@1
^X1o1JeRqfl4ig9KkB1qU:AH;3]HRF76dkc]S2M?6nAW_mpXnOcZYpLR2UTf4`LS
C92A8<]E_<G7X_X5lQpKf<66OYQYa?o<TU^oX`cIOfXHCe2qNWN1dM<;KbNDV@UT
OnVg>\614SYIc<Iq3T0Qg277\o<2<T0@CKh[jU7n`9J>UU8^80EoUTQbbU[U]epm
H6IT?T?2Rp;:R4MfnRD=jS3]EH=UXDcAD5W2k[R:?CEEe@3:\Kh7EcdSQSNTE5[O
hCX`MdY\4OG6pkZA^6e2V1nZHZ2i7X2O5gB40CYbD09`RB3qRGJ=2GV4FTo`IAjT
QX>NFQp7cANgKlIPPq@mLeA1DFUT6DZ1a@l<i[]N3>E?K\aU_pC;6mQ7Zo[gGo88
:CkdR_TYmFh>L4pe;h_QfR<bGq4@\c::q[c3lT8TNmW>MfAb^QBW041_UcW2O@iM
p6VDdXGOHW28Wh`H^B5:G4XEXha^;qZW47IKbG8V6k7_k7FF[Z^6UY]:IUCUGpoM
?aQ`7UZW0FKWI`dK6@U[PRZFGECEk0^L5JeA`l:\gHDQ7qFBe@PbRi5]GlOQb4FQ
c4QYnh2eH_NTY5_?6gjPHK[TX;piR76LSJDlJpKjJ]M6nD[A;3O\D8QK`1R5P_7E
oRkdH;CfO2UVT\4`FcTYgeSNbM5]Q<o5B0nOgIZoeq1bH^<3KR@=9SW\WYhCjYch
qFFTG7f1aI2qF=lIe=N]X@c4C\E=@^?UOLiI8bkBC8oO=O9WBPI1bidAbXY3Z9o5
YfA6VQ9Pk<jQFYUIq<NBk8\`cn0OG^oNbIC]?^UiPjoXn_CKqRQ@O<BNB\iiI9n^
i8i1_RFnef6UCqOgOa]TYP@j9SelH><HTnJXX`?dCp70ZagE]RYmqh;mLLTq4GBc
;b`7g;g<[4SkBHJY6WHg7cZCRVOgqH:NQ>jTdc=Zcj3MKEgXiS<Zqfj1j?BIZN;;
o0m]gPC2iqC`aIHA;`T0Z[A`dHCWdE:0J5^`dVpT9UODCc:kT^d[B3M0Q];6QYY\
Pmc4_?p^@[k6mP5nIcW2_[S]Z;df<Q9WjEaF_XpEDh?BBI84fd\OVjY[VR2e2jPL
Cq<;4GSm36T]KcaDBXf0>a;`fdi=QW3cCbiQFDIF4GZ6fGGPcF4FgBBPdE[7BNF;
U6fVk^n?3dT]KcaDBXf0>a;`fdi=QW3cCbiQFDIF4GZ6fGGPcF4FgBBPdE[7BNF;
U6fVk^n?3dT]KcaDBXf0>a;`fdi=QW3cCbiQFDIF4GZ6fGGPcF4FgBBPdE[7BNF;
U6f`V^fa8Nj7^iR`_?ZC]Rq=a>ciSSf]ZhYSlUC2^2m3E>RjU7CN=WhCBEHGVlS;
a5_JPG3gG;B99o@lBT`mLMU=h0\WMSk]ZhYSlUC2^2m3E>RjU_W79Po5BE6GVlS;
a5_JPG3gG;B99o@lBT`mLMU=h0\WMSk]ZhYSlUC2^2m3E>RjU7CN=WhCBEHGVlS;
a5_JPG3gG;B99o@lBT`mLMU=C?RWmhFCc\NP6dQ28nmpEBeAVU5;>c<c:B85ChX8
9e86cT9koNA;=Lm@T9\ZGmNU_cmn\P@PZ[C=@PhW?eSJEO<G<YL\Gc<m:k7mTcXL
Dk7gmT_lQcA81Tf>[Z;Y7m`^nNNYc5APfWCo23ZL?eSJE>mGWf5k>c<c:B85ChX8
9e86cT9koNA;=Lm@T9\ZGmNU_cmn\P@PZ[C=@PhW?eSJE>1aJfL9INIde4TS_haZ
LoqJVQj5`A^iH2`6MA_A_dEhk>cc1^F=V8A4^:]?F_FnjECCX^Na0f?HRoMe2D0M
=2;=FkHW0A]iH2`6MA_A_dEhk>cc1^F=V8A4^:]?F_FnjECCX^Na0f?HRoMe2D0M
=2;=FkHW0A]iH2`6MA_A_dEhk>cc1^F=V8A4^:]?F_FnjECCX^Na0f?HRoMe2D0M
=2;=fU5]JcWeoXbm8ZFPOkiqMiB4SNKKdl5gFe@pgmkS3mmg3W2m_?e0YL@jUWb_
\475>8gVH6FN861I23Ie0AfepTFgfAmqbW`a@H^?DfTno[lgeK_19CX7[U6FpLmX
Vjf9P3f80L^Q7ZeqDjFTH\gQqWaV]0C_T]W0i3m\6lnIYqNOEQ_c8cj63W6nL@pQ
YO;<V1L7ec@K;oPNmR1pJOV77_LUp<7Mm75955XYVX2kGVN2D]bg?_Pe3GF@_7dK
:n[K7]_dM:3R\C:@ed<X=lPep@oaE:XEg1VqQ7?dKZ\L8^2P@CQ4CZF74Bb[jDIE
QaefQ8WVpcI?[fopSXKS4]b[Jgl_KCNkUU0cWoTq\8IHeOSmXgZUkCadSPmnkH\3
coNkJ[`EU^`qGXO7?o7WP]@WU`cl@AHEYbD]HB5KY3O:;V<Lp6FF2B<F8fSEB8bD
4F]l^]6F;NLSB]UZ]nOA8q_iX7nMhWHdM0cJALZCmPWV:;V>ZeIdJ0[R5ap:aDHV
nkkG5Zb@0LS97EVL[jVEEVAoG<4XRl74`HJD_GeoY1C04WU\o8[q49B2A@ALpYIF
PF0>hTag@8F@8GO^]DVP_\Noj;;bioH3qU_Xh_<nU0ZfEK;kFg7O:fKHHE8=jh?k
\M?I:qZcf8I6hc;KDAUfCafh>hlXV7UF]TB^k]AhNZpAPdf1MU^<BLM^PC?DnSe8
k1G7:bHf0aKgNmFqP]n_7P6bqB[a=I]@KR6ObDgoiD[=@jPH0Na;HFAMj\aUpkZ1
6KYiKJgJgjhmhJXF5UUgn>Eo5X;8W3^aKpQ;XLPdC1d1?ObaFGER3EJKIgje2[WL
2L8bji59q_VEW9oDe6b1]=1[6[h@<o\n]9oF1C^e[fnHNp63fB@Em39WINN1m9gT
C;?J9NOV82P]5Z^UMTqD_jdUh9]p_BdDE2DZI>qCGTL:`pnZXY<nDDlF@9b^2:=4
DEcIP:khp2MKY@:5R;64?OWHG43dp=lK5m^Ue_>m<kf9V3oR]=F5AMK5^gkMXX7U
n3?1DnW6p`XOQ7aLS_lC9n7@lSYeGfBE`RIT?nLmlo9cW_i3LGeVI^MhqC8Pk;d0
S2?JDCF4SR^QMpO?flXeInSBM6gB3Io`;V]8KaFlUfGJSCCR^CbD`6P`Q[LAD?`Q
gXMQ]Ydc>U^RF^mmGU;lW=_0[;Wb=iAJVbM>G<lN>Qg3Y3;ah`JPoX?;DW^d_RM7
ZpMCVmCPmRp>oKhA1DXG8lgPQ`_5S4]@MW^49V?h[ac`9XlW7leSBPDinAZ9[:aq
GPZgB\M2qh`fDPG@p2mR3EXq?_mO3?1:nI_;GkG;?Z4oURNLDVGZNYNA7e2cSGSB
0d8Wchln;Tkc9Vea<kmA6>pf9`2>K>flEV8meN0TGOF=j]Rmhj>4S2gEVe<_U9Xc
2bQZ^<8pj;T>F6i0Em3B[9Z5NZ8I[0QLKFk@5QnjgdZ0BoRmD;^\Ao?jB[;Ok9[k
l6MT55pA;;Lm@?ZDKmED_[kaeBBeY<I7^OCZGnJ1DGYaJ^[?Df<AbfG?X4cAdBK6
NNb>Jp]eSXdV;7<lpY2g;eJpLiQlEj3SZ\D64ZSbD09D1fnGSef3jinU9n0TpY23
MRh4pf^TT=GL3N28AE5\H5EZYH6TX0>Z3Ba4h>ccG=CGjqGH?MnI>c8?0<5_YLAc
;@F7CcDHTB<W5BIOj?_3=@Nbai@h7:;ni3k8:<7EAJe?J7n0i^Ok9M<Ql8MkZU?\
_?lI]LJ>C@l4=`48kH`;]J5eWpYC^QSK0oV;ANRAPmNgBNi6bRTlJYk2mjUmgG=8
JoLnih;D_XCK_b]D<Y=SU23@il3O`@LeI7J`Y\]94m0o4J=LXOh3:KqkFeXPKGBo
n8i<F@BSELcCFL;SL1n3j8I9IoJAT=KL@kSAk07oP785dQn:DE>30p1_=?;H0MHL
9a;MJR7^19?ofFfS_5^Fd[2E4EknR3>g?7k6FegDU59[Mo2`:LAAn8Af[=6RaDB^
fTDiaF;[<YL>5dAdYHqa:2N0kefmBB7XCJ\MY@041M`=GVSjiPCYRC0l3V[G205M
fn`m1a0O@MTFdX;1OH5fmFNAGZacAj5hkRFVlWOThg;3UF3p45J59T2XaZjnH1F\
6`;DiKSgXB\31m02o6_Q8HD<3^83\\Vb[NH>fLgCh8R2j2fi4XP>Z>JGPc8^n=DP
_OHUTQ_PAWCpb>Qd\\YTX27jf1Qf?a;:3eMINh?g3LjjZ@Z593C>C[ZCJdQa^H=J
?jcb0Cc:>WiGbf[PHodRfE3_3_NdUB<n9DOQ4E:p?Y2:Kc>oh7Mam8HSPjmBgm2[
XdoR:KIhfHC3=aJ5LERD_aO<dJDAZ>Y6]b3N7gN\?1G>UjB@[;1T9I0hhZF12oO]
Njmp3U?FJB?aS>Rd=]HFaabk7UfTm4co;Bf_OkO>c@h5jdkiS>UJTm>oBAB@Rcqh
V0KI]3LhTe<ZDCN5T\^`4bV<j4BF6W3@ab`4GL0OP9\LAdE6h\R=P?77Q[4N=pU8
Qje3f^fc8?iiDc5klH@PY?3EN@jke]EZ\LMa>E_R]g8N^LL?jBMWOV?GGHOQq4W1
8AAbGS\CK=J3gb8gofR^T\7JK^2?a;jIT6m5DcM5@nPPmBLCS43pD]kdYnABoI`0
:@A_>cKb5klJfRTXXG1H<GmBm>l1Gb66c5dB0D=o=e\NBHj]p[PI5a500CCLKZ3Y
SnZN>0e<XPIm1OY7lMNUE8UcVXnCjX2dPCI@>M_T@f[fqcSPjXPNHDMQHU:gmbAU
UBQd8A`FnP]f8R3<Rd81GJ;n:A<E`Y0f2@<jQ0f>q[`K_LdlZ23\?0e[_=fD1YHA
\eVSY?FAc4F;5`2O4QLg_3HChXNB<e@YU=oiq72;T6_bXVXPTcdI09QU;F4A=kDQ
P0C]Q[S=UMKUm1ZJZK_5\M7q>>i0^I@i0F98?lKp[1d86P\RMc;Cb\8O@J9ZGME0
3M^2AmnR3O8h9I\\hY?EmYGJolY]9KTeF?M_NPG0[2`Ccffn@:oQcTic2AVM>h\<
FKpAV19d638ph9_cX_h;:?FmkHKeASR7ab305dc7DPXUGbkI@VI^U969oCMd:=JH
MYbe5KfE;Y3i0BolOK_[q7MHE;GK^E6pFdcYgO_gp`fLFNe5BW=l3>_P91nWki\h
UVn=\YPmgTEhHo@hfqNQiFkP31:ORJWXD54SE;lY?hKWj]3;N8mWcnkBJnME4BVb
>7>I<[5\8ECADIZ[@M8L4=9Eo\Pl2bo\<=^K_D<m2?OXS34CmflVR=4X_?I[ZhR>
b:p4kh4S2gD2P21A99PX2jCMR<:G^Gh^RoDT5;A15@^86fF_fKIVBZkfJA1XLjVk
C6\4GhXLE6f6iH[WHT^[2B2I^6?oB7[=6pWU]@nb<VA;[n:o:C5;iP3oJ6fm:1GP
iUWV6>ND7Oa7@VD_]6X_SO0\e4G`LPXQ`>W2ee\gZDSb[V>1X?g;QcXZ5naG7eW6
pXDR6lhFJm6dIh2HNXde@G9Nc_GH0oI1:IQ>Z]GaYH1h=b4@iY1VWJHGIh_<3j<E
>XO[3Zbeo`EZCO8<UTdLm]e_A@DK`G@q0>9YBb57e;Jl9`CQ59]YLbV83FB3WGKV
3eG_BF:;YjGA<f[1;bfcY0XT8ciVg:Zq`H\G`O:2Em`eRT8U29B\[o^OnKiW77`L
]_^C?:kR\@<Ih@E8R>VkYWGbGT3bRo_V9MH;E;SfLQ3];I?bCWgakUkYmT9GYW3q
5m<OR]5kOMkd=Yh4f>PeZ7UPP3iMQT67`6ad<@^NH5AMYdH0c3Ab;1da2EF<R>]2
O5LZ06<>>0Xao;dMNVej8VL@D]bhT01p7FZ1WGh8Fa\e7Xm:lC@9_M49Lm:Xn2]4
lQQod]CWce?Q:fXPOAHFJ5S7R:hY?^54I7@Z:2EEomhU22UBdD3[H`>k\_@;BWnp
`5;TK<7Y8Vbn<58?X<1D=6O6F:TfAQ48>H6RDie:W0>2RJbK:;eQ:c]cC]q\6`>U
<_\]35Xi\TlL^\CNeH9gnZ?^WG58T4C?1gDCh7^4o8CfNJk<?AhV3E4=Cpi63gJ8
mVC@G8SkM0\ZB]9iDWn4kNJnk=e??dK?V9R4=e0]20S1L8kI]TK[k2iYpiWDkHLl
V=Z7:ldo7HI8?YfcXhh?f9X]P6[<JRBg9S`mV0N<ed10PIiQgCRDcqOW0NXlX5M9
9D3?MKP\dNn4biCdOE<inT<T3HJE4M63VI;0<;bNm<8Y1nafAq<=f3EHK_]nbine
XA<?h9cW2oBEQ\7X0SYU]JjdeC7;>\^`T?cm916IG@Tlq>3O\o:Wh\Lh<Qco=M@D
SC7H2EVK@kn>EP;4C_n?cliS>m5cc33Eg\]e95D]pAVdec?b7Ei[4CN8SIKdQS`C
M93SLVeOjn2Vk<^_Mka=JMm9A_;7Mlb1?SMfq61OH\2[nQigR;Il<HO41lVlh`3?
iQie6DBi\o48JkBbkJ6id;=pA8VoK<>gfZ?c;3Bp4i44L\nE>GCI=\9UXh3;ha9R
4HMalV3G\^A=ZIgRNDVjGFFNfGJ`j`HIc6ob^jC=LQ^5BblO18RI=He[oRn3Q51n
UT86kMG6_^lpX7=NHXSgpMLjg6Gm`N_qOgMZU0=ap4<bK>L?p:6Z4V]H^N<Z^Nmq
Q5`Bl]Fdcmq]oRl7hq\Efb0\9>JnRbWc2`@9?MkDnq]gT6c4hl0=3DRN9S=mS6I:
Xf9V70<8LZOh[kNaof3Y[aMFgfkf=0:R<>dSkOBNk`_B01J46aED57XQ_?=mS6I:
Xf9V70<8LZOh[kNaof3e>addm3=K>\WJT8m@FRe1ln9\e=heRpj86WZ]6N1cXin7
MghjeFe=]j9ILbZ=TkLCUJF<RL40f;cIkAZCKhRVhYPYJ[bBdjJbl\7oaal2EaS4
gBhjeFe=]j9ILbZ=TkLCUJF<RL4dn]XSRHER>RlI9j8UUo0Y0FWmm<MTaq4K=@FT
@6_]g4^?TQ:C>KcX@;7d@6Pi\NQZ]8>S5?SB[@mLRCLTJib0FnF9UMeBCfQ>InWf
oY@BFndm96aC>dcX@;7d@6Pi\NQZ]8>S5?S1N6\1:6^g1DNhFVmiTAh>3^H5nU18
`p5f\9KF1`0Z8UiX5YEcCXe45=ml`IEdj=cBeY:Oe\@i=nUNe:HR>i7Y]f1Of]JN
A@\nYL`\a_MJ@>T7?bOmfN48V0lE`PEdj=cBeY:Oe\@i=nUNe:H8Y>GaHfWGR78l
?2iDg9TkaL3FE?7XQC:PpGT8TiBCaI7HL9eU<B81gH?OiS77G1nCZ[UZeGE634Hi
F`hl<YKIVSgiFBVlR346WGeb8`m`PBcgIHU3@0i1f;?<\_Z_X`nai0nY0DbnWHgV
K[_UhBi1;SgiFBVlR346WGeb8`B<05lmJ:WOo9Y1fVSjcBUk8>[=H>R9p57Lg4j9
Cjg8bR:C0dS1DI_S[[^?FBFL^FdI:J;?lEWKfN@fV_j]D5f;8_iQGXa8A:GeH6]Z
J[HoJV1I<HS1GI_S[[^?FBFL^FdI:J;?lEWP[eXBBnZeJ\A052A_PEc25\]<FVO?
Xq]eUdc`_QG5LMmX?UNNQkGjJb\Y_Cn?f<T:[VAGZfeN<<=6hG5@>1\bUbq3;`c4
c84HRJ9i_1HNO2q7lE6WbI?b8plQ1CUapEG1`?O7_To?Z@cokqi2E>mYiq]o6l4U
B<DSC:`5CbbO_4W^9VPP`ZJ2qG@Wk;=qTbi7T5f9Y=>YT5B=7Q_67kSj_Jo^g=>g
7dEVf6]3@g2N]S4:LgGka_\?X_b8F3>\QdnHG_0qk2S>\On2MWc7mik][dVILX2:
<FQ^46OXe4`f:Lj6BhXCiiMl:Cdl^g:eDIYIOGSoLEjT4Un1MWc7mik][dVILX2:
<FQ^46OXe4`f:Lj6BhXCiiMl:Cdl^g:eDIof8QWYW4iM2NVoaV4lq6:BfA:hlVPc
FebKS0dB7oJX_0KX=F>=:L`oD>FV>A[7_IFm;g;@^TCh`LOA4l<kdLE4Vo8hUVPc
FebKS0dB7oJX_0KX=F>=:L`oD>I2AQOhjl`BMShg3lCh5LOZjK?hYZn0DeVH:`@7
hp@EeZ<T0IVFTS7I;K<9egb=TiZVfQ:MUcbMkV\j_ho=:dUEc\VFUjR`O7nn6jbX
;J@gd4Qd>RAU33DI;5VLePb=TiZVfQ:MUcbMkV\j_ho=:dU<TMNnco`KjP:9hC=I
k0U`D1VUPV9cBHp`X>Cn?ceD`T90\EFTO<e?N=58VAk\<]HlL:SK\[o8?_lV`gG6
bi_H1BHLMD[O3Gm`OLQO[L``=^c>G4@ldneLN458VAk\<]HlL:SK\[o8?_l_T:f@
JEo_0CAdnTR3eJJ?1jbPdE1`eFQpC]GL8M<h_Io7:iQZOaXXZ6k\4>:<;0^1NU@:
E>?MIL6;=TJBCUho<RNN0f3=IkQcC[Q4H9YO4i3JE1BT`mFeSk<a2T:_D0^\NU@:
E>CeP87YmRacem=\@7Qil>8P35k_^d?n>Lfe4>bcq6=_em3J0=b>8Aoh6UX\Z>d]
egGBf\OGhJEOa3T0V\ZF9_cC2ZW4[YX]M_VB;40SH6TgbgRFW5H:YXOnl6BV2fOK
^@XhEPYG3<EKNPJH0dj8c>:0;]T]>;i@f8T7AhO_cmOQ4nPb[56ampQ1`QYcBD^5
K1^ffaB`jDHG0YGTYe1jWlHU?G:Z>UDADYPBHm_ToZL9D7?XaEZN;Jq;P_b>Z106
\Q@7]YBdLa6XhggT7_]foER`X^KOEMe9802ZY8D7[LIn4;7^C59TE0e;FgMHdF2d
VC\cU5ZT7];4EJUWmM7K8^j`F9AY0GRhFg3^BQXZUm0g5ikik_TRB8<KE2WfHYUd
F2Jp\dYG\oB`0LJZ5:gDZBP1>EM2O\QiIC>lGEnAMl@<I<5Mo25Y=lFQ;W5cEolU
E<n_\cWGkgi]XO1[T:Mkbdbm49[eo^GH^C>lGEnA?e8^cgc67k1lY7[b\<W>E55Q
?Mgm5g0K>BJjXZ_WpFh5CjfXGHkiPmh7_]6g9]`n:2=9\n4\NhUeb]i[Y]LGj4`o
TUmC90c;XQBO``;<RFZ`M=Nb8Sj9?lm8B>[m>1h<OFi9^n4\NhUeb]i;cknkWi;m
c[cHFGDeK`g<OOU7J0Uj43>3?S\?epLggoN2>0=TKe;;nbnbK85j?LWKH>:S]eEE
CcZ`AG_7;@^06J[VoB;[l:@WK=3_c;Ll`[n03_CegQYe^2VV@Q@1EZnKH6:S]eEE
CcZ`AG_WFTa=NaK`]li]Ld=9PN<HLei8miEJULCnUDqPo;cnk?3lI:>GkB^j7Y5h
ZC\Z;ZnqXoZOZCTTdCI`EKOaEkD?1L0QF2ik1`:_eKM6IdCLFl;L>Jk376RK;CUF
1H;L6hBbXQKY1>>bb\59;7a`l6hQ^R6WF2ik1`:_eKM6IdCLFl42ga>fca6lb[T<
2<oBUQ^\_JSE>Z^\bQ82qFG6JAe`nK?mTdW[l12R\5jUb10X9bNBd@K]]m0m>OW[
>_NOILZ5Cg35<JbT5L`8LFl28nXgB>2A?CS4JlGoNIEU?10X9bNBd@K]]m0m>OW[
>_HA>RYLUPYH1j;IkjiZEBacFlQ_0>NHip2=CLZ1CR=GCWRP5nF[6lHDd;XVoCE`
;?djkaBebKOeZJi=a?Ne<48Y2B:[DhBd3M2A:=D7NZaJTmY^^hX5jGaDd[XVoCE`
;?djkaBebKOeZJi?^bQIEFo76HoQL0ZPJG^e?:7a>kafc8qZ7\54n8U;IOKhd>]o
C``MU\YDilQOMm5@UO`^3cfeGf^EF@B1>S4L7GJdmn7KV0]Zk[Pl7Q>0Gb[W@a\E
:`PMU\YDilQOMm5@UO`^3cfeGf^EF@BjND\[XbcnAhjPchQ4a@P=B2a0QSgqZ6c;
1cn]G\\Rc=<P<WHW7Q>]RX^ESL=^\ZYGL3?P\:Y=?D1QW>I?l`UIfQVN?[>8Z9il
YOmYJmLO:@^jFBHB7Q>]RX^ESL=^\ZYGL3?P\:bWmD1d^A7C9U\6>Ej>m?8Cfnen
jA`;Je90q1AKFWXEW?O\KIIb_fGE^CMllOI<NCo2O3=lSg;WaYCjLP_CBR\c;jkg
g<X\2f7IjSbd]J49MBo^Wm^;6<`AACMllOI<NCo2O3=lSg;Wa<EoeZE<kR5S;o\S
260@HPbkUnc<CfF^?BME5p2BQ9k:9?<WKf5@CJ<nmKcW5bW>>>O16m:MD8d\Io_N
@6lCDCbh^gEn4Nb>9hh]@cHa8SlFQFW5KSaH=dZJ?A8M5\gi>nO16m:MOPUbV@9[
bK^G@QC>FeAn?1d8_]jQU?affTmncZWhhCphH3NbPgc5>kim:BWcXl3N^=HECUi1
K>0LS:@Vh]oE_3:Ofcmd27IL:cdgY=\oSMnHX`lLT]V4VF]B205e8A[9K;lFTXGG
K>]3oBOVF<hA^cjmn1bc`T\JQ>g[Y<XlU8YGSHE\X?U42I@pbHVCN[iR5S]hH69D
E^aFIRLD54hjhP\[2l0HSDJR89Q4WGeJKPTeC@K@2<qZ=Cf?laJ1kA>5ZSMU756Q
R>]6GTK5N:H?4ZALmo<B\EERmiiI3SQ=ekc3Ql[TFn0?J0ndN4_GgaLc4GefmJQD
R>N6GfKhN:R?4ZALm1EG;^:9o_`BTEV:Vjnh60]PHg<OgnIe^L@^@A^pU<jMfJ`h
f8B0I1H9Ug2Z;GF=D?MbS:Sc_d;k`=\;Ye4fmCiMbnS=1M>T?];AH>]b0an7CX`M
7bMGOY_gOSYF]GFFD?MbS:Sc_d;k`=\;M7H_?\ijbnA=`0TFB]L`E^=O\=73\jnM
giOQpXgcIkkYeY;WYBhi6EjM[IN`LDXg6cN5Q4I]7C^FXIcNkA1@H5;MhmW;bJIg
\\gfl27Xf5eVm61bZUak=iYMLI1?8DXg6cm21RjcnKg\[V3l5bL=WBSnhCjY]RT<
eHU_Ce2[j6=j4La=Kp?hIaY1lLkUR[Se^XKLdQ2CEU5BEAaX1k8P1eMYBkj?U[3Q
keMcEUEBCD5PcZl1b8Rk2eFJ4P5aHI0:hMKLdQ2CBNPj2naX1k8PnE9:ZS;W6J3Q
keJ9Hlb_^\TYD27ji6C^i_0`W@ii[ip`NgcEgBFWb0TC2C>bnek\KFOQ^Jo@:iWG
]c`hc`i=Ncn>a^fkeZiZT<A3L=UZ8Ya<FhaI\ZJjA@Kl4K^bnek\KFOQDVoHjWSk
jc7hc`iFbJQIY^3kcnQ>]`Mi0?jW>Hchh<;SFlncNKLqmV=j7>4ECn8YMm21@MNE
CnF>a>B7?:8WMmMcb7fkB\\NW0F]3lbfGF3;>WVR_X[7Ud\KfARJVF5GXfDB@MNE
CnF>a><j8<jlXdji_gJ5D_JFKTWM@=_nmBa>3HNi;H>WAF_B\aAm9h=:qOGIcFLP
F=iD]>Z:?if=IH8T3<1EL3XfaZ?poQ]a[2EX4==<b2_BLA9aAYmec`hd;EEiZ7?Q
`hFZe4k?;`f09Cm5fAN1Fi1>8@f<@MOM3J6L0;ZChe]ILA8UaS>55Sh;;7nklZ?H
2<5ZhbIB;`f0h4mgPE0Bh4Aikg_fM=ET@kD?0l9]q8^I5YCgKlXhFC2^JINAh]Oi
I?HlNe\In@R]jDZFciUD2^<cgBgYiQm@`VLQE3nYYK]LckKcF]S1HLDni9I2V5OD
N?HlNe\In@9_;DZFca9GDPbWU_>YUQ@;1V4`MV666h^?SJU`<j89Tq_D\_MTIa?=
`ogTT;<45o\5Q?W35@<`oje0QlFULmZM]GA?\KEk[gcYfnQU1gMjK@TcbHcVUK]g
;\=WT50QbC`P4PhQb`KlR<F0Q5FU5Mjm0\:89C\[9lU?7NZ3F@:5aS8YDKHk9WKE
f;qXKhf^kF:Xdj@j`jNgS6750PeM;n50Ygi56TR>l?BRQ6eoJQfC?FJ7oC>?YCNL
C?2FGEAHk:C]Xnlj6:0gS<Aj49_AI2dKYgi56TR>cPeY:VgoJQfC7KKjLMkIoQGj
f50`fYN6OIJ]Kccq`H=VcFU\:Ul^G5Kj?Nccj<W_TePbddHTA=l5T:4fdYYIee]C
7WNn8B_B69?3F?XaLGUTD1_5;2N=GTbD?Nccj<W_TjP^hdHRA=l5T:4fdc3Vj`C8
DRAZ2K_hN3?0jdE]eV^L9`QZWUM5q[SP5RC5<Kn=VVNb3AV7`kR5_a:B=_61M;Rb
jVf0mP7@S0gcWaU[Sa1phm:obOgZ0NNQ34\_ES6SMU_:A:=C8949<fCT:XSLJ9h4
GXmkVnPXP6JJ;?;3gMYHV91DXP;e76SJ@4DYES6SMU_:AXT@Rc^OJbC0UXhXFd8o
NeICi[_<CKDhO@b:6U]7b81ia>OD7d7;pV?fA3IKGCc^dbUWGS=S33[Vb;Qmb9e]
`_R@677e?^nGFkPQFmMC]S1LJ_o`T@TRd\>Hl>fKUC[6iC_OhS=S33[Vb;Qmb94Q
>a6]H[XomM7S;hI>?i50W[E[bb3\[TP`TVBB;X;icTjn>pJiYNaXX@WJTH<TWkZ;
EOR290?[?m64AIQ=9^F9T;S4U3XMC]I;GBE]?W7njhN;d0:\dJ6:81PSQXbNlUZ;
ZOT>:X8e?L64AIQ=9^FU6FCEU6C7IFfN=lcjTPFeLc]G_GLhha3IEcg6f@pO:N4\
jnY?_NT9mlB?D2@gg1AObm]cgam>OkW5F]QN820S:>=HEi\0od2hF6m4O5\>d>fb
6o`G=DOA3N>TD2\gXEW9X8K[gam>OkW5nhjI829S:jhHEC\=MWbi5U3LbBbO>f;L
1A7UH3cpnYd6@JIh[3X566HBYYhhJ?9m\3l778diMR?Ymhc@Lh7Ll9YaQ?M^h6jX
5^i]VD>:8l;gKHT5m1_mjQlV`A6[NJeodL^=78diMR?Ymhc@Lh7Ll99aX?k@Aekj
I6Tk<X:Sab>l2_@md;cCpR0<eK06Gi7UmO<G^RR=]iN7V95a[Pjnd8CF]FAldFY5
@FY^36a<6MMa?3<<8<Fi`SDB`5I\omPDX=9GcRRb7HNDJ8ja[Pjnd8CF]FAldFY5
@F_ooad<D3JJhKZI1P<LSDZB<Mg0`dEZ`q9Nj7ZamD5_A;53Z6HZ_79\;cK^nGaQ
eaNYM6UY`bJ]XJC3\;iREYNPCSEME[_B@:95``k=@\RVP=SGho\>J[o\;7K^nGaQ
eaNYM6UY`bJ]XJneN_5JIJ8BLBcPQkO>o2RQ`;ECikR`1JpFDP`WQR7EDeG9?TPm
_V`Y6LlO5<]d>\c6o]`=DYA3NJlD2:Ng1bJbm]a1<>L8k4_nh\fPb:l;Pj]11Kko
d^PF6L;O5<]d>\c6o]`=DYA3N:lhn_oX7nhgZVADfNJIZg6gnSb<;F^;O?jq_^31
4l8iiVQfP7^4dE\hGdUoI7LP3E]dGlTRN`R3DV;QXAfojJm];0LUaG[3q_7Cj@jI
^cV?7g;H=LMi^e;HdJ>QQAbfOKK]_ZiTo=i8ddaEhOl41IT:i=>PSc?1G_=^D1<l
Gc38\___4aYGj=TH9J>QQAbfOKK]_ZiTo=iR7lm^jA:4RCe18]68>iKZAmeZ6M=S
nWf@_p:5^cJWM0ei`[D5FRa]6P[VoBcCU;egVhOV;OFIDo_S]]YATYS3GA:kb:_1
<Imb84K>S;P519WaSA]3699e;jMTY[cCU;egVhOV;OFIDo\03ACoKY;;nbnbK85j
UVjEb6hVAUZ\0=ZO40qLRZgCF:MFbGFklko0=IEglF8X>]0ml?QjWJfe`N4_J<ah
2gn=jdYUN8JKkj0Aol;LcNe]QLjA]lbW]N<6<RQRd0c]D]Rml?QjWJfe`N4\jdRm
3D\3gXQ^jQYNW>kkNLFMG\;gZ`>\F^6pAI_SXf`PP2QahTk53<lckLO>lEKZloC[
?YCNLC?2FGEAH=7[g:Nb2?:^gS6750PeM;b58?ZdIMRO=]?\RQ6eoJQfC?FJ7oC>
?YCNL^fJX=@UCmF<XdbJW_]6a4g6o@IG7m9j8:JX55MHqU>Tg[Mn=Nok6oOS[;j2
ihEHHFX^l:Fj:4P:UTJI>Km>2ofF8^KJ>MTD=>EVBXjKA=DBY`=OUC@8Eg65<k:X
KMJbhgAOJTdPa4P[O4DPeNR3DGSM\3BHaB4\E3XXdbodO?kc:5O<EOAOkq^^bN`E
>4dbAfL4i2HcmFGG`:TeQAcJH1C;[:Xh:8nHe0fRd`1DSeHj1a9edY99HacJ03n@
Gag=2;_]D6Ua_Vdg3I_=eCWa05]U]b@5A3@]gj7W93R;e1m9mPH^VH40NBo_Ui\X
g383anph0;boO_hR7DGZVKef=oEI_U79C;TT5daTAol7IE9c1EaUe]Q@a6PL:`g6
<MDSBH\01AnXPS0IDVJDbjOaI34ZoTM_;a>TUVNTAhF:I;4gOF\IB3fOdAN9<Tgi
_1nNgo1@7Wa:gAe@cbTq]n41ZCR]^\I3VJjML^@d^^OX0o3i9_^1>iDPl[\na1fF
bBhq3kO?gmYo\A:UGkM3[NX9eH^]:M:^H46HDhY9g@PBLnOXc43mSE@co`\R=NYd
_1VEF9Y?5>J0YkK;9:@o^1n_foGV:lScJ46DA5\YOHHPYghYV;T<jJnii=X;E_9D
92FAh4>bf?D=5hUPpDhl9PO;c[mWjJJIbZ\6E;Wg4:n`gS>I4PRY53;A1aRPLJaG
Pj8mokno;CF\NAlUZY5J@Y^Q?aL2YjJEIEOk>JWgO=Q2@SQD0EjYJLiYEJINQ8DX
<Pcm^3Rj^<KC2`5ok4lSHcE`>dbERpBXE?U_n`b1\Ec2Xi=?FdPFBgkc_1L>l6NE
M`ghllk]d>lQ[IC<Lm00>Rf]nQj:[<B3oRi83meSiZ<fBo3l;BDBTPng>[L>l6Hi
^ogkF`9mTg5Q9I<b?8UY^NKhRZKnNYm?AWHkfje3ReqV`SU<e@6DVYXbV70<\`S0
a>]kCnBj[Y6nl?E=nbK>cUSLH0iXn9\KZmE5M[Z:A2QViCnD>@?LUB5`ogWO0]DI
@e3k]F:G0]:;ih3MjQoI3Z`11=0_W?i5\=fiM2:ICIVW`[QR5R1Y^92q7C[U?2q]
GmFD99D^hIW`SWcLOQnK=\de\UiPJ6EXC`TAO@XfE1jW0c67A=>gObGq=TjLnB1L
]jSM?l0S`Y^49^5dgDFif]<DWaNANU31jamZdSdI`U0TUnTd0la@SSGfQ[bL3Y2k
d<M6UHWe=6pgTAdo^ldK0RhH5<580^UB5?H:WiB>Ceed7KU0UIVEgH?k=bbf6=L3
<:2MDQPUO>YaWcACCUm`i^FANZ3KYpT4QOCT3dk<1ZUELn@m0@`G`D8ILc[>7Wmc
fVgBPhM^?6MiaZN\1?kcmInh1?B:`JQgi0N\3?O_ZYOdQ\[^p1\;e@BE=[LYRd0a
OLnqgAc59A4pbj41AepR]:\gWN5f2T_QP1QQ^DJLeiU@f=EOPWp_]CX6i[$
`endprotected
endmodule
