module CHIP(
    clk,
    rst_n,

    in_valid_1,
    in_valid_2,
    in_data,

    out_valid,
    number_2,
    number_4,
    number_6
);

input clk; 
input rst_n;
input in_valid_1;
input in_valid_2;
input [14:0]in_data;

output out_valid;
output number_2;
output number_4;
output number_6;

/**/

wire C_clk;
wire BUF_CLK;

wire C_rst_n;

wire C_in_valid_1;
wire C_in_valid_2;
wire [14:0] C_in_data;

wire C_out_valid;
wire C_number_2;
wire C_number_4;
wire C_number_6;

/**/

CNN CNN ( .clk(BUF_CLK),
	      .rst_n(C_rst_n),
	      .in_valid_1(C_in_valid_1),
	      .in_valid_2(C_in_valid_2),
	      .in_data(C_in_data),
	      .out_valid(C_out_valid),
	      .number_2(C_number_2),
	      .number_4(C_number_4),
	      .number_6(C_number_6));

/**/

CLKBUFX20 buf0 (.Y(BUF_CLK), .A(C_clk));

P8C I_CLK     (.Y(C_clk),        .PU(1'b1),.PD(1'b0),.P(clk),        .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b1),.CEN(1'b0),.A(1'b0));
P8C I_RESET   (.Y(C_rst_n),      .PU(1'b1),.PD(1'b0),.P(rst_n),      .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));

P4C I_VALID_1 (.Y(C_in_valid_1), .PU(1'b1),.PD(1'b0),.P(in_valid_1), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_VALID_2 (.Y(C_in_valid_2), .PU(1'b1),.PD(1'b0),.P(in_valid_2), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));

P4C I_IN_0    (.Y(C_in_data[0]), .PU(1'b1),.PD(1'b0),.P(in_data[0]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_1    (.Y(C_in_data[1]), .PU(1'b1),.PD(1'b0),.P(in_data[1]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_2    (.Y(C_in_data[2]), .PU(1'b1),.PD(1'b0),.P(in_data[2]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_3    (.Y(C_in_data[3]), .PU(1'b1),.PD(1'b0),.P(in_data[3]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_4    (.Y(C_in_data[4]), .PU(1'b1),.PD(1'b0),.P(in_data[4]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_5    (.Y(C_in_data[5]), .PU(1'b1),.PD(1'b0),.P(in_data[5]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_6    (.Y(C_in_data[6]), .PU(1'b1),.PD(1'b0),.P(in_data[6]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_7    (.Y(C_in_data[7]), .PU(1'b1),.PD(1'b0),.P(in_data[7]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_8    (.Y(C_in_data[8]), .PU(1'b1),.PD(1'b0),.P(in_data[8]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_9    (.Y(C_in_data[9]), .PU(1'b1),.PD(1'b0),.P(in_data[9]), .ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_10   (.Y(C_in_data[10]),.PU(1'b1),.PD(1'b0),.P(in_data[10]),.ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_11   (.Y(C_in_data[11]),.PU(1'b1),.PD(1'b0),.P(in_data[11]),.ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_12   (.Y(C_in_data[12]),.PU(1'b1),.PD(1'b0),.P(in_data[12]),.ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_13   (.Y(C_in_data[13]),.PU(1'b1),.PD(1'b0),.P(in_data[13]),.ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));
P4C I_IN_14   (.Y(C_in_data[14]),.PU(1'b1),.PD(1'b0),.P(in_data[14]),.ODEN(1'b0),.OCEN(1'b0),.CSEN(1'b0),.CEN(1'b1),.A(1'b0));

P8C O_VALID   (.PU(1'b1),.PD(1'b0),.P(out_valid),.ODEN(1'b1),.OCEN(1'b1),.CSEN(1'b0),.CEN(1'b1),.A(C_out_valid));

P8C O_NUM_2   (.PU(1'b1),.PD(1'b0),.P(number_2), .ODEN(1'b1),.OCEN(1'b1),.CSEN(1'b0),.CEN(1'b1),.A(C_number_2));
P8C O_NUM_4   (.PU(1'b1),.PD(1'b0),.P(number_4), .ODEN(1'b1),.OCEN(1'b1),.CSEN(1'b0),.CEN(1'b1),.A(C_number_4));
P8C O_NUM_6   (.PU(1'b1),.PD(1'b0),.P(number_6), .ODEN(1'b1),.OCEN(1'b1),.CSEN(1'b0),.CEN(1'b1),.A(C_number_6));

PVDDR VDDP0 ();
PVSSR GNDP0 ();
PVDDR VDDP1 ();
PVSSR GNDP1 ();
PVDDR VDDP2 ();
PVSSR GNDP2 ();
PVDDR VDDP3 ();
PVSSR GNDP3 ();

PVDDC VDDC0 ();
PVSSC GNDC0 ();
PVDDC VDDC1 ();
PVSSC GNDC1 ();
PVDDC VDDC2 ();
PVSSC GNDC2 ();
PVDDC VDDC3 ();
PVSSC GNDC3 ();

endmodule/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : K-2015.06-SP1
// Date      : Tue Jan 16 10:26:09 2018
/////////////////////////////////////////////////////////////


module CNN ( clk, rst_n, in_valid_1, in_valid_2, in_data, out_valid, number_2, 
        number_4, number_6 );
  input [14:0] in_data;
  input clk, rst_n, in_valid_1, in_valid_2;
  output out_valid, number_2, number_4, number_6;
  wire   N17494, N17495, N17496, N17497, N17498, N17499, N17500, N17501,
         N17502, N17503, N17504, N17505, N17506, N17507, N17508, N17509,
         N17510, N17511, N17512, N17513, N17514, N17515, N17516, N17517,
         N17518, N17519, N17520, N17521, N17522, N17523, N17524, N17525,
         N17526, N17527, N17528, N17529, N17530, N17531, N17532, N17533,
         N17534, N17535, N17536, N17537, N17538, N17539, N17540, N17541,
         N17542, N17543, N17544, N17545, N17546, N17547, N17548, N17549,
         N17550, N17551, N17552, N17553, N17554, N17555, N17556, N17557,
         N17631, N17708, N17785, N18014, N18471, N29216, N29217, N29218,
         N29219, N29220, N29221, N29222, N29223, N29224, N29225, N29226,
         N29227, N29228, N29229, N29230, N29231, N29232, N29233, N29234,
         N29235, N29236, N29237, N29238, N29239, N29240, N29241, N29242,
         N29243, N29244, N29245, N29246, N29247, N29248, N29249, N29250,
         N29251, N29252, N29253, N29254, N29255, N29256, N29257, N29258,
         N29259, N29260, N29261, N29262, N29263, N29264, N29265, N29266,
         N29267, N29268, N29269, N29270, N29271, N29272, N29273, N29274,
         N29275, N29276, N29277, N29278, N29279, N29280, N29281, N29282,
         N29283, N29284, N29285, N29286, N29287, N29288, N29289, N29290,
         N29291, N29292, N29293, N29294, N29295, N29296, N29297, N29298,
         N29299, N29300, N29301, N29302, N29303, N29304, N29305, N29306,
         N29307, N29308, N29309, N29310, N29311, N29312, N29313, N29314,
         N29315, N29316, N29317, N29318, N29319, N29320, N29321, N29322,
         N29323, N29324, N29325, N29326, N29327, N29328, N29329, N29330,
         N29331, N29332, N29333, N29334, N29335, N29336, N29337, N29338,
         N29339, N29340, N29341, N29342, N29343, N29344, N29345, N29346,
         N29347, N29348, N29349, N29350, N29496, N29497, N29498, N29499,
         N29500, N30140, N30141, N30142, N30143, N30144, N30145, add_x_358_n5,
         add_x_358_n4, add_x_358_n3, add_x_358_n2, add_x_358_n1, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16636, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         intadd_0_B_2_, intadd_0_B_1_, intadd_0_B_0_, intadd_0_CI,
         intadd_0_SUM_2_, intadd_0_SUM_1_, intadd_0_SUM_0_, intadd_0_n3,
         intadd_0_n2, intadd_0_n1, intadd_1_B_2_, intadd_1_B_1_, intadd_1_B_0_,
         intadd_1_CI, intadd_1_SUM_2_, intadd_1_SUM_1_, intadd_1_SUM_0_,
         intadd_1_n3, intadd_1_n2, intadd_1_n1, intadd_2_B_2_, intadd_2_B_1_,
         intadd_2_B_0_, intadd_2_CI, intadd_2_SUM_2_, intadd_2_SUM_1_,
         intadd_2_SUM_0_, intadd_2_n3, intadd_2_n2, intadd_2_n1,
         DP_OP_5171J1_127_4278_n107, DP_OP_5171J1_127_4278_n101,
         DP_OP_5171J1_127_4278_n98, DP_OP_5171J1_127_4278_n97,
         DP_OP_5171J1_127_4278_n96, DP_OP_5171J1_127_4278_n95,
         DP_OP_5171J1_127_4278_n94, DP_OP_5171J1_127_4278_n93,
         DP_OP_5171J1_127_4278_n91, DP_OP_5171J1_127_4278_n90,
         DP_OP_5171J1_127_4278_n89, DP_OP_5171J1_127_4278_n88,
         DP_OP_5171J1_127_4278_n87, DP_OP_5171J1_127_4278_n86,
         DP_OP_5171J1_127_4278_n85, DP_OP_5171J1_127_4278_n84,
         DP_OP_5171J1_127_4278_n83, DP_OP_5171J1_127_4278_n82,
         DP_OP_5171J1_127_4278_n81, DP_OP_5171J1_127_4278_n76,
         DP_OP_5171J1_127_4278_n67, DP_OP_5171J1_127_4278_n64,
         DP_OP_5171J1_127_4278_n63, DP_OP_5171J1_127_4278_n62,
         DP_OP_5171J1_127_4278_n61, DP_OP_5171J1_127_4278_n60,
         DP_OP_5171J1_127_4278_n59, DP_OP_5171J1_127_4278_n58,
         DP_OP_5171J1_127_4278_n57, DP_OP_5171J1_127_4278_n56,
         DP_OP_5171J1_127_4278_n55, DP_OP_5171J1_127_4278_n54,
         DP_OP_5171J1_127_4278_n53, DP_OP_5171J1_127_4278_n52,
         DP_OP_5171J1_127_4278_n51, DP_OP_5171J1_127_4278_n50,
         DP_OP_5171J1_127_4278_n49, DP_OP_5171J1_127_4278_n48,
         DP_OP_5171J1_127_4278_n47, DP_OP_5171J1_127_4278_n46,
         DP_OP_5171J1_127_4278_n45, DP_OP_5171J1_127_4278_n44,
         DP_OP_5171J1_127_4278_n43, DP_OP_5171J1_127_4278_n42,
         DP_OP_5171J1_127_4278_n41, DP_OP_5171J1_127_4278_n40,
         DP_OP_5171J1_127_4278_n39, DP_OP_5171J1_127_4278_n38,
         DP_OP_5171J1_127_4278_n37, DP_OP_5171J1_127_4278_n36,
         DP_OP_5171J1_127_4278_n35, DP_OP_5171J1_127_4278_n34,
         DP_OP_5171J1_127_4278_n33, DP_OP_5171J1_127_4278_n32,
         DP_OP_5171J1_127_4278_n31, DP_OP_5171J1_127_4278_n29,
         DP_OP_5171J1_127_4278_n28, DP_OP_5171J1_127_4278_n27,
         DP_OP_5171J1_127_4278_n26, DP_OP_5171J1_127_4278_n25,
         DP_OP_5171J1_127_4278_n24, DP_OP_5170J1_126_4278_n107,
         DP_OP_5170J1_126_4278_n101, DP_OP_5170J1_126_4278_n98,
         DP_OP_5170J1_126_4278_n97, DP_OP_5170J1_126_4278_n96,
         DP_OP_5170J1_126_4278_n95, DP_OP_5170J1_126_4278_n94,
         DP_OP_5170J1_126_4278_n93, DP_OP_5170J1_126_4278_n91,
         DP_OP_5170J1_126_4278_n90, DP_OP_5170J1_126_4278_n89,
         DP_OP_5170J1_126_4278_n88, DP_OP_5170J1_126_4278_n87,
         DP_OP_5170J1_126_4278_n86, DP_OP_5170J1_126_4278_n85,
         DP_OP_5170J1_126_4278_n84, DP_OP_5170J1_126_4278_n83,
         DP_OP_5170J1_126_4278_n82, DP_OP_5170J1_126_4278_n81,
         DP_OP_5170J1_126_4278_n76, DP_OP_5170J1_126_4278_n67,
         DP_OP_5170J1_126_4278_n64, DP_OP_5170J1_126_4278_n63,
         DP_OP_5170J1_126_4278_n62, DP_OP_5170J1_126_4278_n61,
         DP_OP_5170J1_126_4278_n60, DP_OP_5170J1_126_4278_n59,
         DP_OP_5170J1_126_4278_n58, DP_OP_5170J1_126_4278_n57,
         DP_OP_5170J1_126_4278_n56, DP_OP_5170J1_126_4278_n55,
         DP_OP_5170J1_126_4278_n54, DP_OP_5170J1_126_4278_n53,
         DP_OP_5170J1_126_4278_n52, DP_OP_5170J1_126_4278_n51,
         DP_OP_5170J1_126_4278_n50, DP_OP_5170J1_126_4278_n49,
         DP_OP_5170J1_126_4278_n48, DP_OP_5170J1_126_4278_n47,
         DP_OP_5170J1_126_4278_n46, DP_OP_5170J1_126_4278_n45,
         DP_OP_5170J1_126_4278_n44, DP_OP_5170J1_126_4278_n43,
         DP_OP_5170J1_126_4278_n42, DP_OP_5170J1_126_4278_n41,
         DP_OP_5170J1_126_4278_n40, DP_OP_5170J1_126_4278_n39,
         DP_OP_5170J1_126_4278_n38, DP_OP_5170J1_126_4278_n37,
         DP_OP_5170J1_126_4278_n36, DP_OP_5170J1_126_4278_n35,
         DP_OP_5170J1_126_4278_n34, DP_OP_5170J1_126_4278_n33,
         DP_OP_5170J1_126_4278_n32, DP_OP_5170J1_126_4278_n31,
         DP_OP_5170J1_126_4278_n29, DP_OP_5170J1_126_4278_n28,
         DP_OP_5170J1_126_4278_n27, DP_OP_5170J1_126_4278_n26,
         DP_OP_5170J1_126_4278_n25, DP_OP_5170J1_126_4278_n24,
         DP_OP_5169J1_125_4278_n107, DP_OP_5169J1_125_4278_n101,
         DP_OP_5169J1_125_4278_n98, DP_OP_5169J1_125_4278_n97,
         DP_OP_5169J1_125_4278_n96, DP_OP_5169J1_125_4278_n95,
         DP_OP_5169J1_125_4278_n94, DP_OP_5169J1_125_4278_n93,
         DP_OP_5169J1_125_4278_n91, DP_OP_5169J1_125_4278_n90,
         DP_OP_5169J1_125_4278_n89, DP_OP_5169J1_125_4278_n88,
         DP_OP_5169J1_125_4278_n87, DP_OP_5169J1_125_4278_n86,
         DP_OP_5169J1_125_4278_n85, DP_OP_5169J1_125_4278_n84,
         DP_OP_5169J1_125_4278_n83, DP_OP_5169J1_125_4278_n82,
         DP_OP_5169J1_125_4278_n81, DP_OP_5169J1_125_4278_n76,
         DP_OP_5169J1_125_4278_n67, DP_OP_5169J1_125_4278_n64,
         DP_OP_5169J1_125_4278_n63, DP_OP_5169J1_125_4278_n62,
         DP_OP_5169J1_125_4278_n61, DP_OP_5169J1_125_4278_n60,
         DP_OP_5169J1_125_4278_n59, DP_OP_5169J1_125_4278_n58,
         DP_OP_5169J1_125_4278_n57, DP_OP_5169J1_125_4278_n56,
         DP_OP_5169J1_125_4278_n55, DP_OP_5169J1_125_4278_n54,
         DP_OP_5169J1_125_4278_n53, DP_OP_5169J1_125_4278_n52,
         DP_OP_5169J1_125_4278_n51, DP_OP_5169J1_125_4278_n50,
         DP_OP_5169J1_125_4278_n49, DP_OP_5169J1_125_4278_n48,
         DP_OP_5169J1_125_4278_n47, DP_OP_5169J1_125_4278_n46,
         DP_OP_5169J1_125_4278_n45, DP_OP_5169J1_125_4278_n44,
         DP_OP_5169J1_125_4278_n43, DP_OP_5169J1_125_4278_n42,
         DP_OP_5169J1_125_4278_n41, DP_OP_5169J1_125_4278_n40,
         DP_OP_5169J1_125_4278_n39, DP_OP_5169J1_125_4278_n38,
         DP_OP_5169J1_125_4278_n37, DP_OP_5169J1_125_4278_n36,
         DP_OP_5169J1_125_4278_n35, DP_OP_5169J1_125_4278_n34,
         DP_OP_5169J1_125_4278_n33, DP_OP_5169J1_125_4278_n32,
         DP_OP_5169J1_125_4278_n31, DP_OP_5169J1_125_4278_n29,
         DP_OP_5169J1_125_4278_n28, DP_OP_5169J1_125_4278_n27,
         DP_OP_5169J1_125_4278_n26, DP_OP_5169J1_125_4278_n25,
         DP_OP_5169J1_125_4278_n24, DP_OP_5168J1_124_9881_n78,
         DP_OP_5168J1_124_9881_n76, DP_OP_5168J1_124_9881_n73,
         DP_OP_5168J1_124_9881_n71, DP_OP_5168J1_124_9881_n70,
         DP_OP_5168J1_124_9881_n67, DP_OP_5168J1_124_9881_n66,
         DP_OP_5168J1_124_9881_n65, DP_OP_5168J1_124_9881_n63,
         DP_OP_5168J1_124_9881_n61, DP_OP_5168J1_124_9881_n60,
         DP_OP_5168J1_124_9881_n58, DP_OP_5168J1_124_9881_n57,
         DP_OP_5168J1_124_9881_n56, DP_OP_5168J1_124_9881_n55,
         DP_OP_5168J1_124_9881_n54, DP_OP_5168J1_124_9881_n53,
         DP_OP_5168J1_124_9881_n48, DP_OP_5168J1_124_9881_n45,
         DP_OP_5168J1_124_9881_n43, DP_OP_5168J1_124_9881_n42,
         DP_OP_5168J1_124_9881_n41, DP_OP_5168J1_124_9881_n40,
         DP_OP_5168J1_124_9881_n39, DP_OP_5168J1_124_9881_n38,
         DP_OP_5168J1_124_9881_n37, DP_OP_5168J1_124_9881_n36,
         DP_OP_5168J1_124_9881_n35, DP_OP_5168J1_124_9881_n34,
         DP_OP_5168J1_124_9881_n33, DP_OP_5168J1_124_9881_n31,
         DP_OP_5168J1_124_9881_n30, DP_OP_5168J1_124_9881_n29,
         DP_OP_5168J1_124_9881_n28, DP_OP_5168J1_124_9881_n27,
         DP_OP_5168J1_124_9881_n26, DP_OP_5168J1_124_9881_n25,
         DP_OP_5168J1_124_9881_n24, DP_OP_5168J1_124_9881_n23,
         DP_OP_5168J1_124_9881_n22, DP_OP_5168J1_124_9881_n21,
         DP_OP_5168J1_124_9881_n20, DP_OP_5168J1_124_9881_n19,
         DP_OP_5168J1_124_9881_n18, DP_OP_5168J1_124_9881_n17,
         DP_OP_5168J1_124_9881_n16, DP_OP_5168J1_124_9881_n15,
         DP_OP_5168J1_124_9881_n14, DP_OP_5168J1_124_9881_n13,
         DP_OP_5168J1_124_9881_n12, DP_OP_5167J1_123_9881_n78,
         DP_OP_5167J1_123_9881_n76, DP_OP_5167J1_123_9881_n73,
         DP_OP_5167J1_123_9881_n71, DP_OP_5167J1_123_9881_n70,
         DP_OP_5167J1_123_9881_n67, DP_OP_5167J1_123_9881_n66,
         DP_OP_5167J1_123_9881_n65, DP_OP_5167J1_123_9881_n63,
         DP_OP_5167J1_123_9881_n61, DP_OP_5167J1_123_9881_n60,
         DP_OP_5167J1_123_9881_n58, DP_OP_5167J1_123_9881_n57,
         DP_OP_5167J1_123_9881_n56, DP_OP_5167J1_123_9881_n55,
         DP_OP_5167J1_123_9881_n54, DP_OP_5167J1_123_9881_n53,
         DP_OP_5167J1_123_9881_n48, DP_OP_5167J1_123_9881_n45,
         DP_OP_5167J1_123_9881_n43, DP_OP_5167J1_123_9881_n42,
         DP_OP_5167J1_123_9881_n41, DP_OP_5167J1_123_9881_n40,
         DP_OP_5167J1_123_9881_n39, DP_OP_5167J1_123_9881_n38,
         DP_OP_5167J1_123_9881_n37, DP_OP_5167J1_123_9881_n36,
         DP_OP_5167J1_123_9881_n35, DP_OP_5167J1_123_9881_n34,
         DP_OP_5167J1_123_9881_n33, DP_OP_5167J1_123_9881_n31,
         DP_OP_5167J1_123_9881_n30, DP_OP_5167J1_123_9881_n29,
         DP_OP_5167J1_123_9881_n28, DP_OP_5167J1_123_9881_n27,
         DP_OP_5167J1_123_9881_n26, DP_OP_5167J1_123_9881_n25,
         DP_OP_5167J1_123_9881_n24, DP_OP_5167J1_123_9881_n23,
         DP_OP_5167J1_123_9881_n22, DP_OP_5167J1_123_9881_n21,
         DP_OP_5167J1_123_9881_n20, DP_OP_5167J1_123_9881_n19,
         DP_OP_5167J1_123_9881_n18, DP_OP_5167J1_123_9881_n17,
         DP_OP_5167J1_123_9881_n16, DP_OP_5167J1_123_9881_n15,
         DP_OP_5167J1_123_9881_n14, DP_OP_5167J1_123_9881_n13,
         DP_OP_5167J1_123_9881_n12, DP_OP_5166J1_122_9881_n78,
         DP_OP_5166J1_122_9881_n76, DP_OP_5166J1_122_9881_n73,
         DP_OP_5166J1_122_9881_n71, DP_OP_5166J1_122_9881_n70,
         DP_OP_5166J1_122_9881_n67, DP_OP_5166J1_122_9881_n66,
         DP_OP_5166J1_122_9881_n65, DP_OP_5166J1_122_9881_n63,
         DP_OP_5166J1_122_9881_n61, DP_OP_5166J1_122_9881_n60,
         DP_OP_5166J1_122_9881_n58, DP_OP_5166J1_122_9881_n57,
         DP_OP_5166J1_122_9881_n56, DP_OP_5166J1_122_9881_n55,
         DP_OP_5166J1_122_9881_n54, DP_OP_5166J1_122_9881_n53,
         DP_OP_5166J1_122_9881_n48, DP_OP_5166J1_122_9881_n45,
         DP_OP_5166J1_122_9881_n43, DP_OP_5166J1_122_9881_n42,
         DP_OP_5166J1_122_9881_n41, DP_OP_5166J1_122_9881_n40,
         DP_OP_5166J1_122_9881_n39, DP_OP_5166J1_122_9881_n38,
         DP_OP_5166J1_122_9881_n37, DP_OP_5166J1_122_9881_n36,
         DP_OP_5166J1_122_9881_n35, DP_OP_5166J1_122_9881_n34,
         DP_OP_5166J1_122_9881_n33, DP_OP_5166J1_122_9881_n31,
         DP_OP_5166J1_122_9881_n30, DP_OP_5166J1_122_9881_n29,
         DP_OP_5166J1_122_9881_n28, DP_OP_5166J1_122_9881_n27,
         DP_OP_5166J1_122_9881_n26, DP_OP_5166J1_122_9881_n25,
         DP_OP_5166J1_122_9881_n24, DP_OP_5166J1_122_9881_n23,
         DP_OP_5166J1_122_9881_n22, DP_OP_5166J1_122_9881_n21,
         DP_OP_5166J1_122_9881_n20, DP_OP_5166J1_122_9881_n19,
         DP_OP_5166J1_122_9881_n18, DP_OP_5166J1_122_9881_n17,
         DP_OP_5166J1_122_9881_n16, DP_OP_5166J1_122_9881_n15,
         DP_OP_5166J1_122_9881_n14, DP_OP_5166J1_122_9881_n13,
         DP_OP_5166J1_122_9881_n12, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
         n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
         n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523,
         n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
         n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
         n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547,
         n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
         n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
         n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
         n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
         n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
         n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
         n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
         n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859,
         n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
         n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
         n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
         n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
         n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931,
         n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
         n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
         n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
         n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
         n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
         n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
         n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
         n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
         n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
         n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
         n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
         n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
         n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
         n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
         n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
         n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
         n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075,
         n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
         n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
         n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
         n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
         n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
         n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147,
         n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
         n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
         n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
         n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
         n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
         n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
         n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315,
         n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
         n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
         n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339,
         n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
         n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363,
         n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
         n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
         n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
         n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
         n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
         n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
         n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
         n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
         n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
         n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467,
         n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
         n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483,
         n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
         n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499,
         n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507,
         n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
         n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
         n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
         n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539,
         n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
         n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555,
         n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
         n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571,
         n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579,
         n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
         n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595,
         n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603,
         n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611,
         n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627,
         n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
         n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643,
         n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651,
         n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
         n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
         n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675,
         n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683,
         n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
         n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699,
         n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
         n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
         n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723,
         n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
         n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
         n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747,
         n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755,
         n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
         n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771,
         n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
         n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787,
         n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795,
         n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
         n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
         n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
         n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827,
         n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
         n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843,
         n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
         n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859,
         n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
         n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
         n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
         n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891,
         n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899,
         n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
         n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915,
         n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
         n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931,
         n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
         n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
         n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
         n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963,
         n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971,
         n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
         n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987,
         n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
         n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003,
         n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
         n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019,
         n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
         n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
         n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043,
         n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
         n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059,
         n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
         n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
         n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083,
         n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091,
         n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
         n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
         n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115,
         n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
         n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131,
         n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
         n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
         n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155,
         n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163,
         n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
         n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
         n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187,
         n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
         n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203,
         n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
         n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
         n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227,
         n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235,
         n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
         n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251,
         n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
         n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
         n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275,
         n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
         n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
         n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299,
         n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
         n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
         n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323,
         n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331,
         n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
         n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
         n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
         n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
         n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371,
         n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
         n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387,
         n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395,
         n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403,
         n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
         n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419,
         n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
         n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
         n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443,
         n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
         n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
         n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467,
         n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475,
         n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
         n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491,
         n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
         n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507,
         n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515,
         n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
         n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
         n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539,
         n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
         n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
         n31556, n31557, n31558, n31560, n31561, n31562, n31563, n31564,
         n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572,
         n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
         n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588,
         n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596,
         n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604,
         n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612,
         n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620,
         n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628,
         n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
         n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644,
         n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
         n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660,
         n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668,
         n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676,
         n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684,
         n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692,
         n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
         n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
         n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716,
         n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
         n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732,
         n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740,
         n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748,
         n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
         n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764,
         n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772,
         n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780,
         n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788,
         n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796,
         n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804,
         n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812,
         n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820,
         n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828,
         n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836,
         n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844,
         n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852,
         n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860,
         n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868,
         n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876,
         n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884,
         n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892,
         n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900,
         n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908,
         n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916,
         n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924,
         n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932,
         n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
         n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948,
         n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956,
         n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964,
         n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972,
         n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980,
         n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988,
         n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996,
         n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004,
         n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012,
         n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
         n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028,
         n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036,
         n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044,
         n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052,
         n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060,
         n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
         n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076,
         n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084,
         n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092,
         n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100,
         n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108,
         n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116,
         n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124,
         n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132,
         n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140,
         n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148,
         n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156,
         n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164,
         n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172,
         n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180,
         n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
         n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196,
         n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204,
         n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212,
         n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220,
         n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228,
         n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236,
         n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244,
         n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252,
         n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260,
         n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268,
         n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276,
         n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
         n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292,
         n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300,
         n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
         n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316,
         n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324,
         n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332,
         n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340,
         n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348,
         n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
         n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364,
         n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372,
         n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380,
         n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388,
         n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396,
         n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404,
         n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412,
         n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420,
         n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428,
         n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436,
         n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444,
         n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452,
         n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460,
         n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468,
         n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476,
         n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484,
         n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492,
         n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500,
         n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508,
         n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516,
         n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524,
         n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532,
         n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540,
         n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548,
         n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556,
         n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
         n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572,
         n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580,
         n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588,
         n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596,
         n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604,
         n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612,
         n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620,
         n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628,
         n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636,
         n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644,
         n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652,
         n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660,
         n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668,
         n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676,
         n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684,
         n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692,
         n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700,
         n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708,
         n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716,
         n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724,
         n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732,
         n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740,
         n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748,
         n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756,
         n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764,
         n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772,
         n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780,
         n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788,
         n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796,
         n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804,
         n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812,
         n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820,
         n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828,
         n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836,
         n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844,
         n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852,
         n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860,
         n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868,
         n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876,
         n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884,
         n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892,
         n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900,
         n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908,
         n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916,
         n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924,
         n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932,
         n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940,
         n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
         n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956,
         n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964,
         n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972,
         n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980,
         n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988,
         n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996,
         n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004,
         n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012,
         n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020,
         n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028,
         n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036,
         n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044,
         n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052,
         n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
         n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068,
         n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076,
         n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084,
         n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092,
         n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100,
         n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108,
         n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116,
         n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124,
         n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132,
         n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140,
         n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148,
         n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156,
         n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164,
         n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
         n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180,
         n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188,
         n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196,
         n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204,
         n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212,
         n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220,
         n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
         n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
         n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244,
         n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252,
         n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260,
         n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
         n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276,
         n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284,
         n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
         n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300,
         n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308,
         n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316,
         n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324,
         n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332,
         n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
         n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348,
         n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
         n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
         n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372,
         n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
         n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388,
         n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396,
         n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
         n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412,
         n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420,
         n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428,
         n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
         n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444,
         n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
         n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460,
         n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468,
         n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476,
         n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484,
         n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492,
         n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500,
         n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508,
         n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516,
         n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
         n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532,
         n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540,
         n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548,
         n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556,
         n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564,
         n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572,
         n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580,
         n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588,
         n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596,
         n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604,
         n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612,
         n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620,
         n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628,
         n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636,
         n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644,
         n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652,
         n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660,
         n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668,
         n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676,
         n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684,
         n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692,
         n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700,
         n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708,
         n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716,
         n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724,
         n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732,
         n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740,
         n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748,
         n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756,
         n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764,
         n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772,
         n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780,
         n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788,
         n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796,
         n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804,
         n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812,
         n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820,
         n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828,
         n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836,
         n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844,
         n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852,
         n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860,
         n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868,
         n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876,
         n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884,
         n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892,
         n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900,
         n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908,
         n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916,
         n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924,
         n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932,
         n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940,
         n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948,
         n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956,
         n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964,
         n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972,
         n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980,
         n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988,
         n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996,
         n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004,
         n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012,
         n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020,
         n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028,
         n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036,
         n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044,
         n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052,
         n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060,
         n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068,
         n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076,
         n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084,
         n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092,
         n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100,
         n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108,
         n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116,
         n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124,
         n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132,
         n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140,
         n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148,
         n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156,
         n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164,
         n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172,
         n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180,
         n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188,
         n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196,
         n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204,
         n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212,
         n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220,
         n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228,
         n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236,
         n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244,
         n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252,
         n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260,
         n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268,
         n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276,
         n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284,
         n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292,
         n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300,
         n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308,
         n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316,
         n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324,
         n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332,
         n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340,
         n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348,
         n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356,
         n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364,
         n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
         n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380,
         n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388,
         n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396,
         n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404,
         n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412,
         n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420,
         n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428,
         n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436,
         n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444,
         n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452,
         n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460,
         n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468,
         n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476,
         n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484,
         n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492,
         n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500,
         n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508,
         n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516,
         n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524,
         n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532,
         n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540,
         n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548,
         n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556,
         n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564,
         n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572,
         n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580,
         n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588,
         n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596,
         n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604,
         n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612,
         n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620,
         n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628,
         n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636,
         n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644,
         n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652,
         n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660,
         n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668,
         n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
         n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684,
         n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692,
         n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700,
         n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708,
         n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716,
         n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724,
         n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732,
         n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740,
         n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748,
         n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756,
         n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764,
         n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772,
         n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780,
         n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788,
         n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796,
         n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804,
         n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812,
         n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820,
         n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828,
         n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836,
         n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844,
         n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852,
         n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860,
         n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868,
         n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876,
         n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884,
         n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892,
         n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900,
         n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908,
         n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916,
         n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924,
         n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932,
         n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940,
         n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948,
         n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956,
         n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964,
         n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972,
         n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980,
         n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988,
         n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996,
         n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004,
         n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012,
         n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020,
         n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028,
         n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036,
         n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044,
         n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052,
         n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060,
         n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068,
         n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076,
         n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084,
         n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092,
         n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100,
         n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108,
         n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116,
         n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124,
         n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132,
         n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140,
         n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148,
         n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156,
         n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164,
         n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172,
         n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180,
         n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188,
         n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196,
         n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204,
         n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212,
         n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220,
         n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228,
         n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236,
         n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244,
         n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252,
         n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260,
         n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268,
         n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276,
         n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284,
         n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292,
         n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300,
         n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308,
         n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316,
         n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324,
         n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332,
         n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340,
         n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348,
         n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356,
         n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364,
         n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372,
         n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380,
         n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388,
         n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396,
         n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404,
         n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412,
         n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420,
         n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428,
         n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436,
         n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444,
         n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452,
         n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460,
         n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468,
         n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476,
         n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484,
         n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492,
         n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500,
         n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508,
         n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516,
         n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524,
         n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532,
         n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540,
         n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548,
         n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556,
         n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564,
         n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572,
         n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580,
         n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588,
         n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596,
         n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604,
         n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612,
         n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620,
         n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628,
         n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636,
         n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644,
         n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652,
         n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660,
         n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668,
         n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676,
         n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684,
         n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692,
         n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700,
         n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708,
         n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716,
         n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724,
         n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732,
         n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740,
         n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748,
         n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756,
         n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764,
         n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772,
         n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780,
         n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788,
         n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796,
         n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804,
         n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812,
         n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820,
         n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828,
         n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836,
         n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844,
         n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852,
         n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860,
         n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868,
         n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876,
         n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884,
         n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892,
         n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900,
         n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908,
         n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916,
         n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924,
         n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932,
         n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940,
         n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948,
         n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956,
         n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964,
         n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972,
         n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980,
         n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988,
         n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996,
         n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004,
         n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012,
         n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020,
         n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028,
         n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036,
         n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044,
         n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052,
         n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060,
         n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068,
         n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076,
         n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084,
         n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092,
         n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100,
         n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108,
         n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116,
         n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124,
         n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132,
         n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140,
         n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148,
         n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156,
         n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164,
         n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172,
         n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180,
         n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188,
         n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196,
         n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204,
         n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212,
         n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220,
         n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228,
         n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236,
         n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244,
         n36245, n36246, n36247, n36248, n36249, n36250,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [53:0] filter_1;
  wire   [53:0] filter_2;
  wire   [53:0] filter_3;
  wire   [5:0] filter_1_bias;
  wire   [5:0] filter_2_bias;
  wire   [5:0] filter_3_bias;
  wire   [2:0] ns;
  wire   [6:0] counter;
  wire   [485:0] weight_1;
  wire   [5:0] weight_1_bias_1;
  wire   [5:0] weight_1_bias_2;
  wire   [5:0] weight_1_bias_3;
  wire   [53:0] weight_2;
  wire   [5:0] weight_2_bias_1;
  wire   [5:0] weight_2_bias_2;
  wire   [5:0] weight_2_bias_3;
  wire   [63:0] pixel;
  wire   [539:0] conv_1;
  wire   [6:5] cursor;
  wire   [539:0] conv_2;
  wire   [539:0] conv_3;
  wire   [134:0] pool;
  wire   [29:0] affine_1;
  wire   [47:0] affine_2;
  wire   [3:0] cs;

  RA1SH R1 ( .Q({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_1}), .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 1'b0}), .CLK(clk), 
        .CEN(1'b0), .OEN(1'b0), .WEN(1'b0) );
  ADDHXL add_x_358_U5 ( .A(n36245), .B(add_x_358_n5), .CO(add_x_358_n4), .S(
        N29497) );
  ADDHXL add_x_358_U4 ( .A(N18014), .B(add_x_358_n4), .CO(add_x_358_n3), .S(
        N29498) );
  ADDHXL add_x_358_U3 ( .A(N18471), .B(add_x_358_n3), .CO(add_x_358_n2), .S(
        N29499) );
  ADDHXL add_x_358_U2 ( .A(n36244), .B(add_x_358_n2), .CO(add_x_358_n1), .S(
        N29500) );
  DFFRHQXL cs_reg_0_ ( .D(ns[0]), .CK(clk), .RN(rst_n), .Q(cs[0]) );
  DFFRHQXL cs_reg_2_ ( .D(ns[2]), .CK(clk), .RN(rst_n), .Q(cs[2]) );
  DFFRHQX2 counter_reg_1_ ( .D(N30140), .CK(clk), .RN(rst_n), .Q(counter[1])
         );
  DFFRHQXL counter_reg_2_ ( .D(N30141), .CK(clk), .RN(rst_n), .Q(counter[2])
         );
  DFFRHQXL counter_reg_4_ ( .D(N30143), .CK(clk), .RN(rst_n), .Q(counter[4])
         );
  DFFRHQXL counter_reg_5_ ( .D(N30144), .CK(clk), .RN(rst_n), .Q(counter[5])
         );
  DFFRHQXL counter_reg_6_ ( .D(N30145), .CK(clk), .RN(rst_n), .Q(counter[6])
         );
  DFFRHQXL cs_reg_1_ ( .D(ns[1]), .CK(clk), .RN(rst_n), .Q(cs[1]) );
  DFFRHQXL pixel_reg_63__0_ ( .D(N17557), .CK(clk), .RN(rst_n), .Q(pixel[63])
         );
  DFFRHQXL pixel_reg_62__0_ ( .D(N17556), .CK(clk), .RN(rst_n), .Q(pixel[62])
         );
  DFFRHQXL pixel_reg_61__0_ ( .D(N17555), .CK(clk), .RN(rst_n), .Q(pixel[61])
         );
  DFFRHQXL pixel_reg_60__0_ ( .D(N17554), .CK(clk), .RN(rst_n), .Q(pixel[60])
         );
  DFFRHQXL pixel_reg_59__0_ ( .D(N17553), .CK(clk), .RN(rst_n), .Q(pixel[59])
         );
  DFFRHQXL pixel_reg_58__0_ ( .D(N17552), .CK(clk), .RN(rst_n), .Q(pixel[58])
         );
  DFFRHQXL pixel_reg_57__0_ ( .D(N17551), .CK(clk), .RN(rst_n), .Q(pixel[57])
         );
  DFFRHQXL pixel_reg_56__0_ ( .D(N17550), .CK(clk), .RN(rst_n), .Q(pixel[56])
         );
  DFFRHQXL pixel_reg_55__0_ ( .D(N17549), .CK(clk), .RN(rst_n), .Q(pixel[55])
         );
  DFFRHQXL pixel_reg_54__0_ ( .D(N17548), .CK(clk), .RN(rst_n), .Q(pixel[54])
         );
  DFFRHQXL pixel_reg_53__0_ ( .D(N17547), .CK(clk), .RN(rst_n), .Q(pixel[53])
         );
  DFFRHQXL pixel_reg_52__0_ ( .D(N17546), .CK(clk), .RN(rst_n), .Q(pixel[52])
         );
  DFFRHQXL pixel_reg_51__0_ ( .D(N17545), .CK(clk), .RN(rst_n), .Q(pixel[51])
         );
  DFFRHQXL pixel_reg_50__0_ ( .D(N17544), .CK(clk), .RN(rst_n), .Q(pixel[50])
         );
  DFFRHQXL pixel_reg_49__0_ ( .D(N17543), .CK(clk), .RN(rst_n), .Q(pixel[49])
         );
  DFFRHQXL pixel_reg_48__0_ ( .D(N17542), .CK(clk), .RN(rst_n), .Q(pixel[48])
         );
  DFFRHQXL pixel_reg_47__0_ ( .D(N17541), .CK(clk), .RN(rst_n), .Q(pixel[47])
         );
  DFFRHQXL pixel_reg_46__0_ ( .D(N17540), .CK(clk), .RN(rst_n), .Q(pixel[46])
         );
  DFFRHQXL pixel_reg_45__0_ ( .D(N17539), .CK(clk), .RN(rst_n), .Q(pixel[45])
         );
  DFFRHQXL pixel_reg_44__0_ ( .D(N17538), .CK(clk), .RN(rst_n), .Q(pixel[44])
         );
  DFFRHQXL pixel_reg_43__0_ ( .D(N17537), .CK(clk), .RN(rst_n), .Q(pixel[43])
         );
  DFFRHQXL pixel_reg_42__0_ ( .D(N17536), .CK(clk), .RN(rst_n), .Q(pixel[42])
         );
  DFFRHQXL pixel_reg_41__0_ ( .D(N17535), .CK(clk), .RN(rst_n), .Q(pixel[41])
         );
  DFFRHQXL pixel_reg_40__0_ ( .D(N17534), .CK(clk), .RN(rst_n), .Q(pixel[40])
         );
  DFFRHQXL pixel_reg_39__0_ ( .D(N17533), .CK(clk), .RN(rst_n), .Q(pixel[39])
         );
  DFFRHQXL pixel_reg_38__0_ ( .D(N17532), .CK(clk), .RN(rst_n), .Q(pixel[38])
         );
  DFFRHQXL pixel_reg_37__0_ ( .D(N17531), .CK(clk), .RN(rst_n), .Q(pixel[37])
         );
  DFFRHQXL pixel_reg_36__0_ ( .D(N17530), .CK(clk), .RN(rst_n), .Q(pixel[36])
         );
  DFFRHQXL pixel_reg_35__0_ ( .D(N17529), .CK(clk), .RN(rst_n), .Q(pixel[35])
         );
  DFFRHQXL pixel_reg_34__0_ ( .D(N17528), .CK(clk), .RN(rst_n), .Q(pixel[34])
         );
  DFFRHQXL pixel_reg_33__0_ ( .D(N17527), .CK(clk), .RN(rst_n), .Q(pixel[33])
         );
  DFFRHQXL pixel_reg_32__0_ ( .D(N17526), .CK(clk), .RN(rst_n), .Q(pixel[32])
         );
  DFFRHQXL pixel_reg_31__0_ ( .D(N17525), .CK(clk), .RN(rst_n), .Q(pixel[31])
         );
  DFFRHQXL pixel_reg_30__0_ ( .D(N17524), .CK(clk), .RN(rst_n), .Q(pixel[30])
         );
  DFFRHQXL pixel_reg_29__0_ ( .D(N17523), .CK(clk), .RN(rst_n), .Q(pixel[29])
         );
  DFFRHQXL pixel_reg_28__0_ ( .D(N17522), .CK(clk), .RN(rst_n), .Q(pixel[28])
         );
  DFFRHQXL pixel_reg_27__0_ ( .D(N17521), .CK(clk), .RN(rst_n), .Q(pixel[27])
         );
  DFFRHQXL pixel_reg_26__0_ ( .D(N17520), .CK(clk), .RN(rst_n), .Q(pixel[26])
         );
  DFFRHQXL pixel_reg_25__0_ ( .D(N17519), .CK(clk), .RN(rst_n), .Q(pixel[25])
         );
  DFFRHQXL pixel_reg_24__0_ ( .D(N17518), .CK(clk), .RN(rst_n), .Q(pixel[24])
         );
  DFFRHQXL pixel_reg_23__0_ ( .D(N17517), .CK(clk), .RN(rst_n), .Q(pixel[23])
         );
  DFFRHQXL pixel_reg_22__0_ ( .D(N17516), .CK(clk), .RN(rst_n), .Q(pixel[22])
         );
  DFFRHQXL pixel_reg_21__0_ ( .D(N17515), .CK(clk), .RN(rst_n), .Q(pixel[21])
         );
  DFFRHQXL pixel_reg_20__0_ ( .D(N17514), .CK(clk), .RN(rst_n), .Q(pixel[20])
         );
  DFFRHQXL pixel_reg_19__0_ ( .D(N17513), .CK(clk), .RN(rst_n), .Q(pixel[19])
         );
  DFFRHQXL pixel_reg_18__0_ ( .D(N17512), .CK(clk), .RN(rst_n), .Q(pixel[18])
         );
  DFFRHQXL pixel_reg_17__0_ ( .D(N17511), .CK(clk), .RN(rst_n), .Q(pixel[17])
         );
  DFFRHQXL pixel_reg_16__0_ ( .D(N17510), .CK(clk), .RN(rst_n), .Q(pixel[16])
         );
  DFFRHQXL pixel_reg_15__0_ ( .D(N17509), .CK(clk), .RN(rst_n), .Q(pixel[15])
         );
  DFFRHQXL pixel_reg_14__0_ ( .D(N17508), .CK(clk), .RN(rst_n), .Q(pixel[14])
         );
  DFFRHQXL pixel_reg_13__0_ ( .D(N17507), .CK(clk), .RN(rst_n), .Q(pixel[13])
         );
  DFFRHQXL pixel_reg_12__0_ ( .D(N17506), .CK(clk), .RN(rst_n), .Q(pixel[12])
         );
  DFFRHQXL pixel_reg_11__0_ ( .D(N17505), .CK(clk), .RN(rst_n), .Q(pixel[11])
         );
  DFFRHQXL pixel_reg_10__0_ ( .D(N17504), .CK(clk), .RN(rst_n), .Q(pixel[10])
         );
  DFFRHQXL pixel_reg_9__0_ ( .D(N17503), .CK(clk), .RN(rst_n), .Q(pixel[9]) );
  DFFRHQXL pixel_reg_8__0_ ( .D(N17502), .CK(clk), .RN(rst_n), .Q(pixel[8]) );
  DFFRHQXL pixel_reg_7__0_ ( .D(N17501), .CK(clk), .RN(rst_n), .Q(pixel[7]) );
  DFFRHQXL pixel_reg_6__0_ ( .D(N17500), .CK(clk), .RN(rst_n), .Q(pixel[6]) );
  DFFRHQXL pixel_reg_5__0_ ( .D(N17499), .CK(clk), .RN(rst_n), .Q(pixel[5]) );
  DFFRHQXL pixel_reg_4__0_ ( .D(N17498), .CK(clk), .RN(rst_n), .Q(pixel[4]) );
  DFFRHQXL pixel_reg_3__0_ ( .D(N17497), .CK(clk), .RN(rst_n), .Q(pixel[3]) );
  DFFRHQXL pixel_reg_2__0_ ( .D(N17496), .CK(clk), .RN(rst_n), .Q(pixel[2]) );
  DFFRHQXL pixel_reg_1__0_ ( .D(N17495), .CK(clk), .RN(rst_n), .Q(pixel[1]) );
  DFFRHQXL pixel_reg_0__0_ ( .D(N17494), .CK(clk), .RN(rst_n), .Q(pixel[0]) );
  DFFRHQX4 cursor_reg_0_ ( .D(n16638), .CK(clk), .RN(rst_n), .Q(N17631) );
  DFFRHQX4 cursor_reg_2_ ( .D(n16640), .CK(clk), .RN(rst_n), .Q(N17785) );
  DFFRHQX4 cursor_reg_4_ ( .D(n16642), .CK(clk), .RN(rst_n), .Q(N18471) );
  DFFRHQXL cursor_reg_6_ ( .D(n16644), .CK(clk), .RN(rst_n), .Q(cursor[6]) );
  DFFRHQXL filter_2_reg_8__5_ ( .D(n14843), .CK(clk), .RN(rst_n), .Q(
        filter_2[53]) );
  DFFRHQXL filter_2_reg_7__5_ ( .D(n14837), .CK(clk), .RN(rst_n), .Q(
        filter_2[47]) );
  DFFRHQXL filter_2_reg_8__4_ ( .D(n14842), .CK(clk), .RN(rst_n), .Q(
        filter_2[52]) );
  DFFRHQXL filter_2_reg_7__4_ ( .D(n14836), .CK(clk), .RN(rst_n), .Q(
        filter_2[46]) );
  DFFRHQXL filter_2_reg_8__3_ ( .D(n14841), .CK(clk), .RN(rst_n), .Q(
        filter_2[51]) );
  DFFRHQXL filter_2_reg_7__3_ ( .D(n14835), .CK(clk), .RN(rst_n), .Q(
        filter_2[45]) );
  DFFRHQXL filter_2_reg_8__2_ ( .D(n14840), .CK(clk), .RN(rst_n), .Q(
        filter_2[50]) );
  DFFRHQXL filter_2_reg_7__2_ ( .D(n14834), .CK(clk), .RN(rst_n), .Q(
        filter_2[44]) );
  DFFRHQXL filter_2_reg_8__1_ ( .D(n14839), .CK(clk), .RN(rst_n), .Q(
        filter_2[49]) );
  DFFRHQXL filter_2_reg_7__1_ ( .D(n14833), .CK(clk), .RN(rst_n), .Q(
        filter_2[43]) );
  DFFRHQXL filter_2_reg_8__0_ ( .D(n14838), .CK(clk), .RN(rst_n), .Q(
        filter_2[48]) );
  DFFRHQXL filter_2_reg_7__0_ ( .D(n14832), .CK(clk), .RN(rst_n), .Q(
        filter_2[42]) );
  DFFRHQXL filter_2_reg_6__5_ ( .D(n14831), .CK(clk), .RN(rst_n), .Q(
        filter_2[41]) );
  DFFRHQXL filter_2_reg_6__4_ ( .D(n14830), .CK(clk), .RN(rst_n), .Q(
        filter_2[40]) );
  DFFRHQXL filter_2_reg_6__3_ ( .D(n14829), .CK(clk), .RN(rst_n), .Q(
        filter_2[39]) );
  DFFRHQXL filter_2_reg_6__2_ ( .D(n14828), .CK(clk), .RN(rst_n), .Q(
        filter_2[38]) );
  DFFRHQXL filter_2_reg_6__1_ ( .D(n14827), .CK(clk), .RN(rst_n), .Q(
        filter_2[37]) );
  DFFRHQXL filter_2_reg_6__0_ ( .D(n14826), .CK(clk), .RN(rst_n), .Q(
        filter_2[36]) );
  DFFRHQXL filter_2_reg_5__5_ ( .D(n14825), .CK(clk), .RN(rst_n), .Q(
        filter_2[35]) );
  DFFRHQXL filter_2_reg_5__4_ ( .D(n14824), .CK(clk), .RN(rst_n), .Q(
        filter_2[34]) );
  DFFRHQXL filter_2_reg_5__3_ ( .D(n14823), .CK(clk), .RN(rst_n), .Q(
        filter_2[33]) );
  DFFRHQXL filter_2_reg_5__2_ ( .D(n14822), .CK(clk), .RN(rst_n), .Q(
        filter_2[32]) );
  DFFRHQXL filter_2_reg_5__1_ ( .D(n14821), .CK(clk), .RN(rst_n), .Q(
        filter_2[31]) );
  DFFRHQXL filter_2_reg_5__0_ ( .D(n14820), .CK(clk), .RN(rst_n), .Q(
        filter_2[30]) );
  DFFRHQXL filter_2_reg_4__5_ ( .D(n14819), .CK(clk), .RN(rst_n), .Q(
        filter_2[29]) );
  DFFRHQXL filter_2_reg_4__4_ ( .D(n14818), .CK(clk), .RN(rst_n), .Q(
        filter_2[28]) );
  DFFRHQXL filter_2_reg_4__3_ ( .D(n14817), .CK(clk), .RN(rst_n), .Q(
        filter_2[27]) );
  DFFRHQXL filter_2_reg_4__2_ ( .D(n14816), .CK(clk), .RN(rst_n), .Q(
        filter_2[26]) );
  DFFRHQXL filter_2_reg_4__1_ ( .D(n14815), .CK(clk), .RN(rst_n), .Q(
        filter_2[25]) );
  DFFRHQXL filter_2_reg_4__0_ ( .D(n14814), .CK(clk), .RN(rst_n), .Q(
        filter_2[24]) );
  DFFRHQXL filter_2_reg_3__5_ ( .D(n14813), .CK(clk), .RN(rst_n), .Q(
        filter_2[23]) );
  DFFRHQXL filter_2_reg_3__4_ ( .D(n14812), .CK(clk), .RN(rst_n), .Q(
        filter_2[22]) );
  DFFRHQXL filter_2_reg_3__3_ ( .D(n14811), .CK(clk), .RN(rst_n), .Q(
        filter_2[21]) );
  DFFRHQXL filter_2_reg_3__2_ ( .D(n14810), .CK(clk), .RN(rst_n), .Q(
        filter_2[20]) );
  DFFRHQXL filter_2_reg_3__1_ ( .D(n14809), .CK(clk), .RN(rst_n), .Q(
        filter_2[19]) );
  DFFRHQXL filter_2_reg_3__0_ ( .D(n14808), .CK(clk), .RN(rst_n), .Q(
        filter_2[18]) );
  DFFRHQXL filter_2_reg_2__5_ ( .D(n14807), .CK(clk), .RN(rst_n), .Q(
        filter_2[17]) );
  DFFRHQXL filter_2_reg_2__4_ ( .D(n14806), .CK(clk), .RN(rst_n), .Q(
        filter_2[16]) );
  DFFRHQXL filter_2_reg_2__3_ ( .D(n14805), .CK(clk), .RN(rst_n), .Q(
        filter_2[15]) );
  DFFRHQXL filter_2_reg_2__2_ ( .D(n14804), .CK(clk), .RN(rst_n), .Q(
        filter_2[14]) );
  DFFRHQXL filter_2_reg_2__1_ ( .D(n14803), .CK(clk), .RN(rst_n), .Q(
        filter_2[13]) );
  DFFRHQXL filter_2_reg_2__0_ ( .D(n14802), .CK(clk), .RN(rst_n), .Q(
        filter_2[12]) );
  DFFRHQXL filter_2_reg_1__5_ ( .D(n14801), .CK(clk), .RN(rst_n), .Q(
        filter_2[11]) );
  DFFRHQXL filter_2_reg_1__4_ ( .D(n14800), .CK(clk), .RN(rst_n), .Q(
        filter_2[10]) );
  DFFRHQXL filter_2_reg_1__3_ ( .D(n14799), .CK(clk), .RN(rst_n), .Q(
        filter_2[9]) );
  DFFRHQXL filter_2_reg_1__2_ ( .D(n14798), .CK(clk), .RN(rst_n), .Q(
        filter_2[8]) );
  DFFRHQXL filter_2_reg_1__1_ ( .D(n14797), .CK(clk), .RN(rst_n), .Q(
        filter_2[7]) );
  DFFRHQXL filter_2_reg_1__0_ ( .D(n14796), .CK(clk), .RN(rst_n), .Q(
        filter_2[6]) );
  DFFRHQXL filter_2_reg_0__0_ ( .D(n14795), .CK(clk), .RN(rst_n), .Q(
        filter_2[0]) );
  DFFRHQXL filter_2_reg_0__5_ ( .D(n14794), .CK(clk), .RN(rst_n), .Q(
        filter_2[5]) );
  DFFRHQXL filter_2_reg_0__4_ ( .D(n14793), .CK(clk), .RN(rst_n), .Q(
        filter_2[4]) );
  DFFRHQXL filter_2_reg_0__3_ ( .D(n14792), .CK(clk), .RN(rst_n), .Q(
        filter_2[3]) );
  DFFRHQXL filter_2_reg_0__2_ ( .D(n14791), .CK(clk), .RN(rst_n), .Q(
        filter_2[2]) );
  DFFRHQXL filter_2_reg_0__1_ ( .D(n14790), .CK(clk), .RN(rst_n), .Q(
        filter_2[1]) );
  DFFRHQXL filter_3_reg_8__5_ ( .D(n14789), .CK(clk), .RN(rst_n), .Q(
        filter_3[53]) );
  DFFRHQXL filter_3_reg_8__4_ ( .D(n14788), .CK(clk), .RN(rst_n), .Q(
        filter_3[52]) );
  DFFRHQXL filter_3_reg_8__3_ ( .D(n14787), .CK(clk), .RN(rst_n), .Q(
        filter_3[51]) );
  DFFRHQXL filter_3_reg_8__2_ ( .D(n14786), .CK(clk), .RN(rst_n), .Q(
        filter_3[50]) );
  DFFRHQXL filter_3_reg_8__1_ ( .D(n14785), .CK(clk), .RN(rst_n), .Q(
        filter_3[49]) );
  DFFRHQXL filter_3_reg_8__0_ ( .D(n14784), .CK(clk), .RN(rst_n), .Q(
        filter_3[48]) );
  DFFRHQXL filter_3_reg_7__5_ ( .D(n14783), .CK(clk), .RN(rst_n), .Q(
        filter_3[47]) );
  DFFRHQXL filter_3_reg_7__4_ ( .D(n14782), .CK(clk), .RN(rst_n), .Q(
        filter_3[46]) );
  DFFRHQXL filter_3_reg_7__3_ ( .D(n14781), .CK(clk), .RN(rst_n), .Q(
        filter_3[45]) );
  DFFRHQXL filter_3_reg_7__2_ ( .D(n14780), .CK(clk), .RN(rst_n), .Q(
        filter_3[44]) );
  DFFRHQXL filter_3_reg_7__1_ ( .D(n14779), .CK(clk), .RN(rst_n), .Q(
        filter_3[43]) );
  DFFRHQXL filter_3_reg_7__0_ ( .D(n14778), .CK(clk), .RN(rst_n), .Q(
        filter_3[42]) );
  DFFRHQXL filter_3_reg_6__5_ ( .D(n14777), .CK(clk), .RN(rst_n), .Q(
        filter_3[41]) );
  DFFRHQXL filter_3_reg_6__4_ ( .D(n14776), .CK(clk), .RN(rst_n), .Q(
        filter_3[40]) );
  DFFRHQXL filter_3_reg_6__3_ ( .D(n14775), .CK(clk), .RN(rst_n), .Q(
        filter_3[39]) );
  DFFRHQXL filter_3_reg_6__2_ ( .D(n14774), .CK(clk), .RN(rst_n), .Q(
        filter_3[38]) );
  DFFRHQXL filter_3_reg_6__1_ ( .D(n14773), .CK(clk), .RN(rst_n), .Q(
        filter_3[37]) );
  DFFRHQXL filter_3_reg_6__0_ ( .D(n14772), .CK(clk), .RN(rst_n), .Q(
        filter_3[36]) );
  DFFRHQXL filter_3_reg_5__5_ ( .D(n14771), .CK(clk), .RN(rst_n), .Q(
        filter_3[35]) );
  DFFRHQXL filter_3_reg_5__4_ ( .D(n14770), .CK(clk), .RN(rst_n), .Q(
        filter_3[34]) );
  DFFRHQXL filter_3_reg_5__3_ ( .D(n14769), .CK(clk), .RN(rst_n), .Q(
        filter_3[33]) );
  DFFRHQXL filter_3_reg_5__2_ ( .D(n14768), .CK(clk), .RN(rst_n), .Q(
        filter_3[32]) );
  DFFRHQXL filter_3_reg_5__1_ ( .D(n14767), .CK(clk), .RN(rst_n), .Q(
        filter_3[31]) );
  DFFRHQXL filter_3_reg_5__0_ ( .D(n14766), .CK(clk), .RN(rst_n), .Q(
        filter_3[30]) );
  DFFRHQXL filter_3_reg_4__5_ ( .D(n14765), .CK(clk), .RN(rst_n), .Q(
        filter_3[29]) );
  DFFRHQXL filter_3_reg_4__4_ ( .D(n14764), .CK(clk), .RN(rst_n), .Q(
        filter_3[28]) );
  DFFRHQXL filter_3_reg_4__3_ ( .D(n14763), .CK(clk), .RN(rst_n), .Q(
        filter_3[27]) );
  DFFRHQXL filter_3_reg_4__2_ ( .D(n14762), .CK(clk), .RN(rst_n), .Q(
        filter_3[26]) );
  DFFRHQXL filter_3_reg_4__1_ ( .D(n14761), .CK(clk), .RN(rst_n), .Q(
        filter_3[25]) );
  DFFRHQXL filter_3_reg_4__0_ ( .D(n14760), .CK(clk), .RN(rst_n), .Q(
        filter_3[24]) );
  DFFRHQXL filter_3_reg_3__5_ ( .D(n14759), .CK(clk), .RN(rst_n), .Q(
        filter_3[23]) );
  DFFRHQXL filter_3_reg_3__4_ ( .D(n14758), .CK(clk), .RN(rst_n), .Q(
        filter_3[22]) );
  DFFRHQXL filter_3_reg_3__3_ ( .D(n14757), .CK(clk), .RN(rst_n), .Q(
        filter_3[21]) );
  DFFRHQXL filter_3_reg_3__2_ ( .D(n14756), .CK(clk), .RN(rst_n), .Q(
        filter_3[20]) );
  DFFRHQXL filter_3_reg_3__1_ ( .D(n14755), .CK(clk), .RN(rst_n), .Q(
        filter_3[19]) );
  DFFRHQXL filter_3_reg_3__0_ ( .D(n14754), .CK(clk), .RN(rst_n), .Q(
        filter_3[18]) );
  DFFRHQXL filter_3_reg_2__5_ ( .D(n14753), .CK(clk), .RN(rst_n), .Q(
        filter_3[17]) );
  DFFRHQXL filter_3_reg_2__4_ ( .D(n14752), .CK(clk), .RN(rst_n), .Q(
        filter_3[16]) );
  DFFRHQXL filter_3_reg_2__3_ ( .D(n14751), .CK(clk), .RN(rst_n), .Q(
        filter_3[15]) );
  DFFRHQXL filter_3_reg_2__2_ ( .D(n14750), .CK(clk), .RN(rst_n), .Q(
        filter_3[14]) );
  DFFRHQXL filter_3_reg_2__1_ ( .D(n14749), .CK(clk), .RN(rst_n), .Q(
        filter_3[13]) );
  DFFRHQXL filter_3_reg_2__0_ ( .D(n14748), .CK(clk), .RN(rst_n), .Q(
        filter_3[12]) );
  DFFRHQXL filter_3_reg_1__5_ ( .D(n14747), .CK(clk), .RN(rst_n), .Q(
        filter_3[11]) );
  DFFRHQXL filter_3_reg_1__4_ ( .D(n14746), .CK(clk), .RN(rst_n), .Q(
        filter_3[10]) );
  DFFRHQXL filter_3_reg_1__3_ ( .D(n14745), .CK(clk), .RN(rst_n), .Q(
        filter_3[9]) );
  DFFRHQXL filter_3_reg_1__2_ ( .D(n14744), .CK(clk), .RN(rst_n), .Q(
        filter_3[8]) );
  DFFRHQXL filter_3_reg_1__1_ ( .D(n14743), .CK(clk), .RN(rst_n), .Q(
        filter_3[7]) );
  DFFRHQXL filter_3_reg_1__0_ ( .D(n14742), .CK(clk), .RN(rst_n), .Q(
        filter_3[6]) );
  DFFRHQXL filter_3_reg_0__0_ ( .D(n14741), .CK(clk), .RN(rst_n), .Q(
        filter_3[0]) );
  DFFRHQXL filter_3_reg_0__5_ ( .D(n14740), .CK(clk), .RN(rst_n), .Q(
        filter_3[5]) );
  DFFRHQXL filter_3_reg_0__4_ ( .D(n14739), .CK(clk), .RN(rst_n), .Q(
        filter_3[4]) );
  DFFRHQXL filter_3_reg_0__3_ ( .D(n14738), .CK(clk), .RN(rst_n), .Q(
        filter_3[3]) );
  DFFRHQXL filter_3_reg_0__2_ ( .D(n14737), .CK(clk), .RN(rst_n), .Q(
        filter_3[2]) );
  DFFRHQXL filter_3_reg_0__1_ ( .D(n14736), .CK(clk), .RN(rst_n), .Q(
        filter_3[1]) );
  DFFRHQXL filter_3_bias_reg_0_ ( .D(n14735), .CK(clk), .RN(rst_n), .Q(
        filter_3_bias[0]) );
  DFFRHQXL filter_2_bias_reg_0_ ( .D(n14734), .CK(clk), .RN(rst_n), .Q(
        filter_2_bias[0]) );
  DFFRHQXL filter_1_bias_reg_0_ ( .D(n14733), .CK(clk), .RN(rst_n), .Q(
        filter_1_bias[0]) );
  DFFRHQXL filter_3_bias_reg_5_ ( .D(n14732), .CK(clk), .RN(rst_n), .Q(
        filter_3_bias[5]) );
  DFFRHQXL conv_3_reg_0__14_ ( .D(n15734), .CK(clk), .RN(rst_n), .Q(conv_3[14]) );
  DFFRHQXL conv_3_reg_0__0_ ( .D(n15923), .CK(clk), .RN(rst_n), .Q(conv_3[0])
         );
  DFFRHQXL conv_3_reg_0__5_ ( .D(n15743), .CK(clk), .RN(rst_n), .Q(conv_3[5])
         );
  DFFRHQXL conv_3_reg_0__6_ ( .D(n15742), .CK(clk), .RN(rst_n), .Q(conv_3[6])
         );
  DFFRHQXL conv_3_reg_0__7_ ( .D(n15741), .CK(clk), .RN(rst_n), .Q(conv_3[7])
         );
  DFFRHQXL conv_3_reg_0__8_ ( .D(n15740), .CK(clk), .RN(rst_n), .Q(conv_3[8])
         );
  DFFRHQXL conv_3_reg_0__9_ ( .D(n15739), .CK(clk), .RN(rst_n), .Q(conv_3[9])
         );
  DFFRHQXL conv_3_reg_0__10_ ( .D(n15738), .CK(clk), .RN(rst_n), .Q(conv_3[10]) );
  DFFRHQXL conv_3_reg_0__11_ ( .D(n15737), .CK(clk), .RN(rst_n), .Q(conv_3[11]) );
  DFFRHQXL conv_3_reg_0__12_ ( .D(n15736), .CK(clk), .RN(rst_n), .Q(conv_3[12]) );
  DFFRHQXL conv_3_reg_0__13_ ( .D(n15735), .CK(clk), .RN(rst_n), .Q(conv_3[13]) );
  DFFRHQXL conv_3_reg_1__14_ ( .D(n15724), .CK(clk), .RN(rst_n), .Q(conv_3[29]) );
  DFFRHQXL conv_3_reg_1__0_ ( .D(n15922), .CK(clk), .RN(rst_n), .Q(conv_3[15])
         );
  DFFRHQXL conv_3_reg_1__5_ ( .D(n15733), .CK(clk), .RN(rst_n), .Q(conv_3[20])
         );
  DFFRHQXL conv_3_reg_1__6_ ( .D(n15732), .CK(clk), .RN(rst_n), .Q(conv_3[21])
         );
  DFFRHQXL conv_3_reg_1__7_ ( .D(n15731), .CK(clk), .RN(rst_n), .Q(conv_3[22])
         );
  DFFRHQXL conv_3_reg_1__8_ ( .D(n15730), .CK(clk), .RN(rst_n), .Q(conv_3[23])
         );
  DFFRHQXL conv_3_reg_1__9_ ( .D(n15729), .CK(clk), .RN(rst_n), .Q(conv_3[24])
         );
  DFFRHQXL conv_3_reg_1__10_ ( .D(n15728), .CK(clk), .RN(rst_n), .Q(conv_3[25]) );
  DFFRHQXL conv_3_reg_1__11_ ( .D(n15727), .CK(clk), .RN(rst_n), .Q(conv_3[26]) );
  DFFRHQXL conv_3_reg_1__12_ ( .D(n15726), .CK(clk), .RN(rst_n), .Q(conv_3[27]) );
  DFFRHQXL conv_3_reg_1__13_ ( .D(n15725), .CK(clk), .RN(rst_n), .Q(conv_3[28]) );
  DFFRHQXL conv_3_reg_2__14_ ( .D(n15714), .CK(clk), .RN(rst_n), .Q(conv_3[44]) );
  DFFRHQXL conv_3_reg_2__0_ ( .D(n15921), .CK(clk), .RN(rst_n), .Q(conv_3[30])
         );
  DFFRHQXL conv_3_reg_2__5_ ( .D(n15723), .CK(clk), .RN(rst_n), .Q(conv_3[35])
         );
  DFFRHQXL conv_3_reg_2__6_ ( .D(n15722), .CK(clk), .RN(rst_n), .Q(conv_3[36])
         );
  DFFRHQXL conv_3_reg_2__7_ ( .D(n15721), .CK(clk), .RN(rst_n), .Q(conv_3[37])
         );
  DFFRHQXL conv_3_reg_2__8_ ( .D(n15720), .CK(clk), .RN(rst_n), .Q(conv_3[38])
         );
  DFFRHQXL conv_3_reg_2__9_ ( .D(n15719), .CK(clk), .RN(rst_n), .Q(conv_3[39])
         );
  DFFRHQXL conv_3_reg_2__10_ ( .D(n15718), .CK(clk), .RN(rst_n), .Q(conv_3[40]) );
  DFFRHQXL conv_3_reg_2__11_ ( .D(n15717), .CK(clk), .RN(rst_n), .Q(conv_3[41]) );
  DFFRHQXL conv_3_reg_2__12_ ( .D(n15716), .CK(clk), .RN(rst_n), .Q(conv_3[42]) );
  DFFRHQXL conv_3_reg_2__13_ ( .D(n15715), .CK(clk), .RN(rst_n), .Q(conv_3[43]) );
  DFFRHQXL conv_3_reg_3__14_ ( .D(n15704), .CK(clk), .RN(rst_n), .Q(conv_3[59]) );
  DFFRHQXL conv_3_reg_3__0_ ( .D(n15920), .CK(clk), .RN(rst_n), .Q(conv_3[45])
         );
  DFFRHQXL conv_3_reg_3__5_ ( .D(n15713), .CK(clk), .RN(rst_n), .Q(conv_3[50])
         );
  DFFRHQXL conv_3_reg_3__6_ ( .D(n15712), .CK(clk), .RN(rst_n), .Q(conv_3[51])
         );
  DFFRHQXL conv_3_reg_3__7_ ( .D(n15711), .CK(clk), .RN(rst_n), .Q(conv_3[52])
         );
  DFFRHQXL conv_3_reg_3__8_ ( .D(n15710), .CK(clk), .RN(rst_n), .Q(conv_3[53])
         );
  DFFRHQXL conv_3_reg_3__9_ ( .D(n15709), .CK(clk), .RN(rst_n), .Q(conv_3[54])
         );
  DFFRHQXL conv_3_reg_3__10_ ( .D(n15708), .CK(clk), .RN(rst_n), .Q(conv_3[55]) );
  DFFRHQXL conv_3_reg_3__11_ ( .D(n15707), .CK(clk), .RN(rst_n), .Q(conv_3[56]) );
  DFFRHQXL conv_3_reg_3__12_ ( .D(n15706), .CK(clk), .RN(rst_n), .Q(conv_3[57]) );
  DFFRHQXL conv_3_reg_3__13_ ( .D(n15705), .CK(clk), .RN(rst_n), .Q(conv_3[58]) );
  DFFRHQXL conv_3_reg_4__14_ ( .D(n15694), .CK(clk), .RN(rst_n), .Q(conv_3[74]) );
  DFFRHQXL conv_3_reg_4__0_ ( .D(n15919), .CK(clk), .RN(rst_n), .Q(conv_3[60])
         );
  DFFRHQXL conv_3_reg_4__5_ ( .D(n15703), .CK(clk), .RN(rst_n), .Q(conv_3[65])
         );
  DFFRHQXL conv_3_reg_4__6_ ( .D(n15702), .CK(clk), .RN(rst_n), .Q(conv_3[66])
         );
  DFFRHQXL conv_3_reg_4__7_ ( .D(n15701), .CK(clk), .RN(rst_n), .Q(conv_3[67])
         );
  DFFRHQXL conv_3_reg_4__8_ ( .D(n15700), .CK(clk), .RN(rst_n), .Q(conv_3[68])
         );
  DFFRHQXL conv_3_reg_4__9_ ( .D(n15699), .CK(clk), .RN(rst_n), .Q(conv_3[69])
         );
  DFFRHQXL conv_3_reg_4__10_ ( .D(n15698), .CK(clk), .RN(rst_n), .Q(conv_3[70]) );
  DFFRHQXL conv_3_reg_4__11_ ( .D(n15697), .CK(clk), .RN(rst_n), .Q(conv_3[71]) );
  DFFRHQXL conv_3_reg_4__12_ ( .D(n15696), .CK(clk), .RN(rst_n), .Q(conv_3[72]) );
  DFFRHQXL conv_3_reg_4__13_ ( .D(n15695), .CK(clk), .RN(rst_n), .Q(conv_3[73]) );
  DFFRHQXL conv_3_reg_5__14_ ( .D(n15684), .CK(clk), .RN(rst_n), .Q(conv_3[89]) );
  DFFRHQXL conv_3_reg_5__0_ ( .D(n15918), .CK(clk), .RN(rst_n), .Q(conv_3[75])
         );
  DFFRHQXL conv_3_reg_5__5_ ( .D(n15693), .CK(clk), .RN(rst_n), .Q(conv_3[80])
         );
  DFFRHQXL conv_3_reg_5__6_ ( .D(n15692), .CK(clk), .RN(rst_n), .Q(conv_3[81])
         );
  DFFRHQXL conv_3_reg_5__7_ ( .D(n15691), .CK(clk), .RN(rst_n), .Q(conv_3[82])
         );
  DFFRHQXL conv_3_reg_5__8_ ( .D(n15690), .CK(clk), .RN(rst_n), .Q(conv_3[83])
         );
  DFFRHQXL conv_3_reg_5__9_ ( .D(n15689), .CK(clk), .RN(rst_n), .Q(conv_3[84])
         );
  DFFRHQXL conv_3_reg_5__10_ ( .D(n15688), .CK(clk), .RN(rst_n), .Q(conv_3[85]) );
  DFFRHQXL conv_3_reg_5__11_ ( .D(n15687), .CK(clk), .RN(rst_n), .Q(conv_3[86]) );
  DFFRHQXL conv_3_reg_5__12_ ( .D(n15686), .CK(clk), .RN(rst_n), .Q(conv_3[87]) );
  DFFRHQXL conv_3_reg_5__13_ ( .D(n15685), .CK(clk), .RN(rst_n), .Q(conv_3[88]) );
  DFFRHQXL conv_3_reg_6__14_ ( .D(n15674), .CK(clk), .RN(rst_n), .Q(
        conv_3[104]) );
  DFFRHQXL conv_3_reg_6__0_ ( .D(n15917), .CK(clk), .RN(rst_n), .Q(conv_3[90])
         );
  DFFRHQXL conv_3_reg_6__5_ ( .D(n15683), .CK(clk), .RN(rst_n), .Q(conv_3[95])
         );
  DFFRHQXL conv_3_reg_6__6_ ( .D(n15682), .CK(clk), .RN(rst_n), .Q(conv_3[96])
         );
  DFFRHQXL conv_3_reg_6__7_ ( .D(n15681), .CK(clk), .RN(rst_n), .Q(conv_3[97])
         );
  DFFRHQXL conv_3_reg_6__8_ ( .D(n15680), .CK(clk), .RN(rst_n), .Q(conv_3[98])
         );
  DFFRHQXL conv_3_reg_6__9_ ( .D(n15679), .CK(clk), .RN(rst_n), .Q(conv_3[99])
         );
  DFFRHQXL conv_3_reg_6__10_ ( .D(n15678), .CK(clk), .RN(rst_n), .Q(
        conv_3[100]) );
  DFFRHQXL conv_3_reg_6__11_ ( .D(n15677), .CK(clk), .RN(rst_n), .Q(
        conv_3[101]) );
  DFFRHQXL conv_3_reg_6__12_ ( .D(n15676), .CK(clk), .RN(rst_n), .Q(
        conv_3[102]) );
  DFFRHQXL conv_3_reg_6__13_ ( .D(n15675), .CK(clk), .RN(rst_n), .Q(
        conv_3[103]) );
  DFFRHQXL conv_3_reg_7__14_ ( .D(n15664), .CK(clk), .RN(rst_n), .Q(
        conv_3[119]) );
  DFFRHQXL conv_3_reg_7__0_ ( .D(n15916), .CK(clk), .RN(rst_n), .Q(conv_3[105]) );
  DFFRHQXL conv_3_reg_7__5_ ( .D(n15673), .CK(clk), .RN(rst_n), .Q(conv_3[110]) );
  DFFRHQXL conv_3_reg_7__6_ ( .D(n15672), .CK(clk), .RN(rst_n), .Q(conv_3[111]) );
  DFFRHQXL conv_3_reg_7__7_ ( .D(n15671), .CK(clk), .RN(rst_n), .Q(conv_3[112]) );
  DFFRHQXL conv_3_reg_7__8_ ( .D(n15670), .CK(clk), .RN(rst_n), .Q(conv_3[113]) );
  DFFRHQXL conv_3_reg_7__9_ ( .D(n15669), .CK(clk), .RN(rst_n), .Q(conv_3[114]) );
  DFFRHQXL conv_3_reg_7__10_ ( .D(n15668), .CK(clk), .RN(rst_n), .Q(
        conv_3[115]) );
  DFFRHQXL conv_3_reg_7__11_ ( .D(n15667), .CK(clk), .RN(rst_n), .Q(
        conv_3[116]) );
  DFFRHQXL conv_3_reg_7__12_ ( .D(n15666), .CK(clk), .RN(rst_n), .Q(
        conv_3[117]) );
  DFFRHQXL conv_3_reg_7__13_ ( .D(n15665), .CK(clk), .RN(rst_n), .Q(
        conv_3[118]) );
  DFFRHQXL conv_3_reg_8__14_ ( .D(n15654), .CK(clk), .RN(rst_n), .Q(
        conv_3[134]) );
  DFFRHQXL conv_3_reg_8__0_ ( .D(n15915), .CK(clk), .RN(rst_n), .Q(conv_3[120]) );
  DFFRHQXL conv_3_reg_8__5_ ( .D(n15663), .CK(clk), .RN(rst_n), .Q(conv_3[125]) );
  DFFRHQXL conv_3_reg_8__6_ ( .D(n15662), .CK(clk), .RN(rst_n), .Q(conv_3[126]) );
  DFFRHQXL conv_3_reg_8__7_ ( .D(n15661), .CK(clk), .RN(rst_n), .Q(conv_3[127]) );
  DFFRHQXL conv_3_reg_8__8_ ( .D(n15660), .CK(clk), .RN(rst_n), .Q(conv_3[128]) );
  DFFRHQXL conv_3_reg_8__9_ ( .D(n15659), .CK(clk), .RN(rst_n), .Q(conv_3[129]) );
  DFFRHQXL conv_3_reg_8__10_ ( .D(n15658), .CK(clk), .RN(rst_n), .Q(
        conv_3[130]) );
  DFFRHQXL conv_3_reg_8__11_ ( .D(n15657), .CK(clk), .RN(rst_n), .Q(
        conv_3[131]) );
  DFFRHQXL conv_3_reg_8__12_ ( .D(n15656), .CK(clk), .RN(rst_n), .Q(
        conv_3[132]) );
  DFFRHQXL conv_3_reg_8__13_ ( .D(n15655), .CK(clk), .RN(rst_n), .Q(
        conv_3[133]) );
  DFFRHQXL conv_3_reg_9__14_ ( .D(n15644), .CK(clk), .RN(rst_n), .Q(
        conv_3[149]) );
  DFFRHQXL conv_3_reg_9__0_ ( .D(n15914), .CK(clk), .RN(rst_n), .Q(conv_3[135]) );
  DFFRHQXL conv_3_reg_9__5_ ( .D(n15653), .CK(clk), .RN(rst_n), .Q(conv_3[140]) );
  DFFRHQXL conv_3_reg_9__6_ ( .D(n15652), .CK(clk), .RN(rst_n), .Q(conv_3[141]) );
  DFFRHQXL conv_3_reg_9__7_ ( .D(n15651), .CK(clk), .RN(rst_n), .Q(conv_3[142]) );
  DFFRHQXL conv_3_reg_9__8_ ( .D(n15650), .CK(clk), .RN(rst_n), .Q(conv_3[143]) );
  DFFRHQXL conv_3_reg_9__9_ ( .D(n15649), .CK(clk), .RN(rst_n), .Q(conv_3[144]) );
  DFFRHQXL conv_3_reg_9__10_ ( .D(n15648), .CK(clk), .RN(rst_n), .Q(
        conv_3[145]) );
  DFFRHQXL conv_3_reg_9__11_ ( .D(n15647), .CK(clk), .RN(rst_n), .Q(
        conv_3[146]) );
  DFFRHQXL conv_3_reg_9__12_ ( .D(n15646), .CK(clk), .RN(rst_n), .Q(
        conv_3[147]) );
  DFFRHQXL conv_3_reg_9__13_ ( .D(n15645), .CK(clk), .RN(rst_n), .Q(
        conv_3[148]) );
  DFFRHQXL conv_3_reg_10__14_ ( .D(n15634), .CK(clk), .RN(rst_n), .Q(
        conv_3[164]) );
  DFFRHQXL conv_3_reg_10__0_ ( .D(n15913), .CK(clk), .RN(rst_n), .Q(
        conv_3[150]) );
  DFFRHQXL conv_3_reg_10__5_ ( .D(n15643), .CK(clk), .RN(rst_n), .Q(
        conv_3[155]) );
  DFFRHQXL conv_3_reg_10__6_ ( .D(n15642), .CK(clk), .RN(rst_n), .Q(
        conv_3[156]) );
  DFFRHQXL conv_3_reg_10__7_ ( .D(n15641), .CK(clk), .RN(rst_n), .Q(
        conv_3[157]) );
  DFFRHQXL conv_3_reg_10__8_ ( .D(n15640), .CK(clk), .RN(rst_n), .Q(
        conv_3[158]) );
  DFFRHQXL conv_3_reg_10__9_ ( .D(n15639), .CK(clk), .RN(rst_n), .Q(
        conv_3[159]) );
  DFFRHQXL conv_3_reg_10__10_ ( .D(n15638), .CK(clk), .RN(rst_n), .Q(
        conv_3[160]) );
  DFFRHQXL conv_3_reg_10__11_ ( .D(n15637), .CK(clk), .RN(rst_n), .Q(
        conv_3[161]) );
  DFFRHQXL conv_3_reg_10__12_ ( .D(n15636), .CK(clk), .RN(rst_n), .Q(
        conv_3[162]) );
  DFFRHQXL conv_3_reg_10__13_ ( .D(n15635), .CK(clk), .RN(rst_n), .Q(
        conv_3[163]) );
  DFFRHQXL conv_3_reg_11__14_ ( .D(n15624), .CK(clk), .RN(rst_n), .Q(
        conv_3[179]) );
  DFFRHQXL conv_3_reg_11__0_ ( .D(n15912), .CK(clk), .RN(rst_n), .Q(
        conv_3[165]) );
  DFFRHQXL conv_3_reg_11__5_ ( .D(n15633), .CK(clk), .RN(rst_n), .Q(
        conv_3[170]) );
  DFFRHQXL conv_3_reg_11__6_ ( .D(n15632), .CK(clk), .RN(rst_n), .Q(
        conv_3[171]) );
  DFFRHQXL conv_3_reg_11__7_ ( .D(n15631), .CK(clk), .RN(rst_n), .Q(
        conv_3[172]) );
  DFFRHQXL conv_3_reg_11__8_ ( .D(n15630), .CK(clk), .RN(rst_n), .Q(
        conv_3[173]) );
  DFFRHQXL conv_3_reg_11__9_ ( .D(n15629), .CK(clk), .RN(rst_n), .Q(
        conv_3[174]) );
  DFFRHQXL conv_3_reg_11__10_ ( .D(n15628), .CK(clk), .RN(rst_n), .Q(
        conv_3[175]) );
  DFFRHQXL conv_3_reg_11__11_ ( .D(n15627), .CK(clk), .RN(rst_n), .Q(
        conv_3[176]) );
  DFFRHQXL conv_3_reg_11__12_ ( .D(n15626), .CK(clk), .RN(rst_n), .Q(
        conv_3[177]) );
  DFFRHQXL conv_3_reg_11__13_ ( .D(n15625), .CK(clk), .RN(rst_n), .Q(
        conv_3[178]) );
  DFFRHQXL conv_3_reg_12__14_ ( .D(n15614), .CK(clk), .RN(rst_n), .Q(
        conv_3[194]) );
  DFFRHQXL conv_3_reg_12__0_ ( .D(n15911), .CK(clk), .RN(rst_n), .Q(
        conv_3[180]) );
  DFFRHQXL conv_3_reg_12__5_ ( .D(n15623), .CK(clk), .RN(rst_n), .Q(
        conv_3[185]) );
  DFFRHQXL conv_3_reg_12__6_ ( .D(n15622), .CK(clk), .RN(rst_n), .Q(
        conv_3[186]) );
  DFFRHQXL conv_3_reg_12__7_ ( .D(n15621), .CK(clk), .RN(rst_n), .Q(
        conv_3[187]) );
  DFFRHQXL conv_3_reg_12__8_ ( .D(n15620), .CK(clk), .RN(rst_n), .Q(
        conv_3[188]) );
  DFFRHQXL conv_3_reg_12__9_ ( .D(n15619), .CK(clk), .RN(rst_n), .Q(
        conv_3[189]) );
  DFFRHQXL conv_3_reg_12__10_ ( .D(n15618), .CK(clk), .RN(rst_n), .Q(
        conv_3[190]) );
  DFFRHQXL conv_3_reg_12__11_ ( .D(n15617), .CK(clk), .RN(rst_n), .Q(
        conv_3[191]) );
  DFFRHQXL conv_3_reg_12__12_ ( .D(n15616), .CK(clk), .RN(rst_n), .Q(
        conv_3[192]) );
  DFFRHQXL conv_3_reg_12__13_ ( .D(n15615), .CK(clk), .RN(rst_n), .Q(
        conv_3[193]) );
  DFFRHQXL conv_3_reg_13__14_ ( .D(n15604), .CK(clk), .RN(rst_n), .Q(
        conv_3[209]) );
  DFFRHQXL conv_3_reg_13__0_ ( .D(n15910), .CK(clk), .RN(rst_n), .Q(
        conv_3[195]) );
  DFFRHQXL conv_3_reg_13__5_ ( .D(n15613), .CK(clk), .RN(rst_n), .Q(
        conv_3[200]) );
  DFFRHQXL conv_3_reg_13__6_ ( .D(n15612), .CK(clk), .RN(rst_n), .Q(
        conv_3[201]) );
  DFFRHQXL conv_3_reg_13__7_ ( .D(n15611), .CK(clk), .RN(rst_n), .Q(
        conv_3[202]) );
  DFFRHQXL conv_3_reg_13__8_ ( .D(n15610), .CK(clk), .RN(rst_n), .Q(
        conv_3[203]) );
  DFFRHQXL conv_3_reg_13__9_ ( .D(n15609), .CK(clk), .RN(rst_n), .Q(
        conv_3[204]) );
  DFFRHQXL conv_3_reg_13__10_ ( .D(n15608), .CK(clk), .RN(rst_n), .Q(
        conv_3[205]) );
  DFFRHQXL conv_3_reg_13__11_ ( .D(n15607), .CK(clk), .RN(rst_n), .Q(
        conv_3[206]) );
  DFFRHQXL conv_3_reg_13__12_ ( .D(n15606), .CK(clk), .RN(rst_n), .Q(
        conv_3[207]) );
  DFFRHQXL conv_3_reg_13__13_ ( .D(n15605), .CK(clk), .RN(rst_n), .Q(
        conv_3[208]) );
  DFFRHQXL conv_3_reg_14__14_ ( .D(n15594), .CK(clk), .RN(rst_n), .Q(
        conv_3[224]) );
  DFFRHQXL conv_3_reg_14__0_ ( .D(n15909), .CK(clk), .RN(rst_n), .Q(
        conv_3[210]) );
  DFFRHQXL conv_3_reg_14__5_ ( .D(n15603), .CK(clk), .RN(rst_n), .Q(
        conv_3[215]) );
  DFFRHQXL conv_3_reg_14__6_ ( .D(n15602), .CK(clk), .RN(rst_n), .Q(
        conv_3[216]) );
  DFFRHQXL conv_3_reg_14__7_ ( .D(n15601), .CK(clk), .RN(rst_n), .Q(
        conv_3[217]) );
  DFFRHQXL conv_3_reg_14__8_ ( .D(n15600), .CK(clk), .RN(rst_n), .Q(
        conv_3[218]) );
  DFFRHQXL conv_3_reg_14__9_ ( .D(n15599), .CK(clk), .RN(rst_n), .Q(
        conv_3[219]) );
  DFFRHQXL conv_3_reg_14__10_ ( .D(n15598), .CK(clk), .RN(rst_n), .Q(
        conv_3[220]) );
  DFFRHQXL conv_3_reg_14__11_ ( .D(n15597), .CK(clk), .RN(rst_n), .Q(
        conv_3[221]) );
  DFFRHQXL conv_3_reg_14__12_ ( .D(n15596), .CK(clk), .RN(rst_n), .Q(
        conv_3[222]) );
  DFFRHQXL conv_3_reg_14__13_ ( .D(n15595), .CK(clk), .RN(rst_n), .Q(
        conv_3[223]) );
  DFFRHQXL conv_3_reg_15__14_ ( .D(n15584), .CK(clk), .RN(rst_n), .Q(
        conv_3[239]) );
  DFFRHQXL conv_3_reg_15__0_ ( .D(n15908), .CK(clk), .RN(rst_n), .Q(
        conv_3[225]) );
  DFFRHQXL conv_3_reg_15__5_ ( .D(n15593), .CK(clk), .RN(rst_n), .Q(
        conv_3[230]) );
  DFFRHQXL conv_3_reg_15__6_ ( .D(n15592), .CK(clk), .RN(rst_n), .Q(
        conv_3[231]) );
  DFFRHQXL conv_3_reg_15__7_ ( .D(n15591), .CK(clk), .RN(rst_n), .Q(
        conv_3[232]) );
  DFFRHQXL conv_3_reg_15__8_ ( .D(n15590), .CK(clk), .RN(rst_n), .Q(
        conv_3[233]) );
  DFFRHQXL conv_3_reg_15__9_ ( .D(n15589), .CK(clk), .RN(rst_n), .Q(
        conv_3[234]) );
  DFFRHQXL conv_3_reg_15__10_ ( .D(n15588), .CK(clk), .RN(rst_n), .Q(
        conv_3[235]) );
  DFFRHQXL conv_3_reg_15__11_ ( .D(n15587), .CK(clk), .RN(rst_n), .Q(
        conv_3[236]) );
  DFFRHQXL conv_3_reg_15__12_ ( .D(n15586), .CK(clk), .RN(rst_n), .Q(
        conv_3[237]) );
  DFFRHQXL conv_3_reg_15__13_ ( .D(n15585), .CK(clk), .RN(rst_n), .Q(
        conv_3[238]) );
  DFFRHQXL conv_3_reg_16__14_ ( .D(n15574), .CK(clk), .RN(rst_n), .Q(
        conv_3[254]) );
  DFFRHQXL conv_3_reg_16__0_ ( .D(n15907), .CK(clk), .RN(rst_n), .Q(
        conv_3[240]) );
  DFFRHQXL conv_3_reg_16__5_ ( .D(n15583), .CK(clk), .RN(rst_n), .Q(
        conv_3[245]) );
  DFFRHQXL conv_3_reg_16__6_ ( .D(n15582), .CK(clk), .RN(rst_n), .Q(
        conv_3[246]) );
  DFFRHQXL conv_3_reg_16__7_ ( .D(n15581), .CK(clk), .RN(rst_n), .Q(
        conv_3[247]) );
  DFFRHQXL conv_3_reg_16__8_ ( .D(n15580), .CK(clk), .RN(rst_n), .Q(
        conv_3[248]) );
  DFFRHQXL conv_3_reg_16__9_ ( .D(n15579), .CK(clk), .RN(rst_n), .Q(
        conv_3[249]) );
  DFFRHQXL conv_3_reg_16__10_ ( .D(n15578), .CK(clk), .RN(rst_n), .Q(
        conv_3[250]) );
  DFFRHQXL conv_3_reg_16__11_ ( .D(n15577), .CK(clk), .RN(rst_n), .Q(
        conv_3[251]) );
  DFFRHQXL conv_3_reg_16__12_ ( .D(n15576), .CK(clk), .RN(rst_n), .Q(
        conv_3[252]) );
  DFFRHQXL conv_3_reg_16__13_ ( .D(n15575), .CK(clk), .RN(rst_n), .Q(
        conv_3[253]) );
  DFFRHQXL conv_3_reg_17__14_ ( .D(n15564), .CK(clk), .RN(rst_n), .Q(
        conv_3[269]) );
  DFFRHQXL conv_3_reg_17__0_ ( .D(n15906), .CK(clk), .RN(rst_n), .Q(
        conv_3[255]) );
  DFFRHQXL conv_3_reg_17__5_ ( .D(n15573), .CK(clk), .RN(rst_n), .Q(
        conv_3[260]) );
  DFFRHQXL conv_3_reg_17__6_ ( .D(n15572), .CK(clk), .RN(rst_n), .Q(
        conv_3[261]) );
  DFFRHQXL conv_3_reg_17__7_ ( .D(n15571), .CK(clk), .RN(rst_n), .Q(
        conv_3[262]) );
  DFFRHQXL conv_3_reg_17__8_ ( .D(n15570), .CK(clk), .RN(rst_n), .Q(
        conv_3[263]) );
  DFFRHQXL conv_3_reg_17__9_ ( .D(n15569), .CK(clk), .RN(rst_n), .Q(
        conv_3[264]) );
  DFFRHQXL conv_3_reg_17__10_ ( .D(n15568), .CK(clk), .RN(rst_n), .Q(
        conv_3[265]) );
  DFFRHQXL conv_3_reg_17__11_ ( .D(n15567), .CK(clk), .RN(rst_n), .Q(
        conv_3[266]) );
  DFFRHQXL conv_3_reg_17__12_ ( .D(n15566), .CK(clk), .RN(rst_n), .Q(
        conv_3[267]) );
  DFFRHQXL conv_3_reg_17__13_ ( .D(n15565), .CK(clk), .RN(rst_n), .Q(
        conv_3[268]) );
  DFFRHQXL conv_3_reg_18__14_ ( .D(n15554), .CK(clk), .RN(rst_n), .Q(
        conv_3[284]) );
  DFFRHQXL conv_3_reg_18__0_ ( .D(n15905), .CK(clk), .RN(rst_n), .Q(
        conv_3[270]) );
  DFFRHQXL conv_3_reg_18__5_ ( .D(n15563), .CK(clk), .RN(rst_n), .Q(
        conv_3[275]) );
  DFFRHQXL conv_3_reg_18__6_ ( .D(n15562), .CK(clk), .RN(rst_n), .Q(
        conv_3[276]) );
  DFFRHQXL conv_3_reg_18__7_ ( .D(n15561), .CK(clk), .RN(rst_n), .Q(
        conv_3[277]) );
  DFFRHQXL conv_3_reg_18__8_ ( .D(n15560), .CK(clk), .RN(rst_n), .Q(
        conv_3[278]) );
  DFFRHQXL conv_3_reg_18__9_ ( .D(n15559), .CK(clk), .RN(rst_n), .Q(
        conv_3[279]) );
  DFFRHQXL conv_3_reg_18__10_ ( .D(n15558), .CK(clk), .RN(rst_n), .Q(
        conv_3[280]) );
  DFFRHQXL conv_3_reg_18__11_ ( .D(n15557), .CK(clk), .RN(rst_n), .Q(
        conv_3[281]) );
  DFFRHQXL conv_3_reg_18__12_ ( .D(n15556), .CK(clk), .RN(rst_n), .Q(
        conv_3[282]) );
  DFFRHQXL conv_3_reg_18__13_ ( .D(n15555), .CK(clk), .RN(rst_n), .Q(
        conv_3[283]) );
  DFFRHQXL conv_3_reg_19__14_ ( .D(n15544), .CK(clk), .RN(rst_n), .Q(
        conv_3[299]) );
  DFFRHQXL conv_3_reg_19__0_ ( .D(n15904), .CK(clk), .RN(rst_n), .Q(
        conv_3[285]) );
  DFFRHQXL conv_3_reg_19__5_ ( .D(n15553), .CK(clk), .RN(rst_n), .Q(
        conv_3[290]) );
  DFFRHQXL conv_3_reg_19__6_ ( .D(n15552), .CK(clk), .RN(rst_n), .Q(
        conv_3[291]) );
  DFFRHQXL conv_3_reg_19__7_ ( .D(n15551), .CK(clk), .RN(rst_n), .Q(
        conv_3[292]) );
  DFFRHQXL conv_3_reg_19__8_ ( .D(n15550), .CK(clk), .RN(rst_n), .Q(
        conv_3[293]) );
  DFFRHQXL conv_3_reg_19__9_ ( .D(n15549), .CK(clk), .RN(rst_n), .Q(
        conv_3[294]) );
  DFFRHQXL conv_3_reg_19__10_ ( .D(n15548), .CK(clk), .RN(rst_n), .Q(
        conv_3[295]) );
  DFFRHQXL conv_3_reg_19__11_ ( .D(n15547), .CK(clk), .RN(rst_n), .Q(
        conv_3[296]) );
  DFFRHQXL conv_3_reg_19__12_ ( .D(n15546), .CK(clk), .RN(rst_n), .Q(
        conv_3[297]) );
  DFFRHQXL conv_3_reg_19__13_ ( .D(n15545), .CK(clk), .RN(rst_n), .Q(
        conv_3[298]) );
  DFFRHQXL conv_3_reg_20__14_ ( .D(n15534), .CK(clk), .RN(rst_n), .Q(
        conv_3[314]) );
  DFFRHQXL conv_3_reg_20__0_ ( .D(n15903), .CK(clk), .RN(rst_n), .Q(
        conv_3[300]) );
  DFFRHQXL conv_3_reg_20__5_ ( .D(n15543), .CK(clk), .RN(rst_n), .Q(
        conv_3[305]) );
  DFFRHQXL conv_3_reg_20__6_ ( .D(n15542), .CK(clk), .RN(rst_n), .Q(
        conv_3[306]) );
  DFFRHQXL conv_3_reg_20__7_ ( .D(n15541), .CK(clk), .RN(rst_n), .Q(
        conv_3[307]) );
  DFFRHQXL conv_3_reg_20__8_ ( .D(n15540), .CK(clk), .RN(rst_n), .Q(
        conv_3[308]) );
  DFFRHQXL conv_3_reg_20__9_ ( .D(n15539), .CK(clk), .RN(rst_n), .Q(
        conv_3[309]) );
  DFFRHQXL conv_3_reg_20__10_ ( .D(n15538), .CK(clk), .RN(rst_n), .Q(
        conv_3[310]) );
  DFFRHQXL conv_3_reg_20__11_ ( .D(n15537), .CK(clk), .RN(rst_n), .Q(
        conv_3[311]) );
  DFFRHQXL conv_3_reg_20__12_ ( .D(n15536), .CK(clk), .RN(rst_n), .Q(
        conv_3[312]) );
  DFFRHQXL conv_3_reg_20__13_ ( .D(n15535), .CK(clk), .RN(rst_n), .Q(
        conv_3[313]) );
  DFFRHQXL conv_3_reg_21__14_ ( .D(n15524), .CK(clk), .RN(rst_n), .Q(
        conv_3[329]) );
  DFFRHQXL conv_3_reg_21__0_ ( .D(n15902), .CK(clk), .RN(rst_n), .Q(
        conv_3[315]) );
  DFFRHQXL conv_3_reg_21__5_ ( .D(n15533), .CK(clk), .RN(rst_n), .Q(
        conv_3[320]) );
  DFFRHQXL conv_3_reg_21__6_ ( .D(n15532), .CK(clk), .RN(rst_n), .Q(
        conv_3[321]) );
  DFFRHQXL conv_3_reg_21__7_ ( .D(n15531), .CK(clk), .RN(rst_n), .Q(
        conv_3[322]) );
  DFFRHQXL conv_3_reg_21__8_ ( .D(n15530), .CK(clk), .RN(rst_n), .Q(
        conv_3[323]) );
  DFFRHQXL conv_3_reg_21__9_ ( .D(n15529), .CK(clk), .RN(rst_n), .Q(
        conv_3[324]) );
  DFFRHQXL conv_3_reg_21__10_ ( .D(n15528), .CK(clk), .RN(rst_n), .Q(
        conv_3[325]) );
  DFFRHQXL conv_3_reg_21__11_ ( .D(n15527), .CK(clk), .RN(rst_n), .Q(
        conv_3[326]) );
  DFFRHQXL conv_3_reg_21__12_ ( .D(n15526), .CK(clk), .RN(rst_n), .Q(
        conv_3[327]) );
  DFFRHQXL conv_3_reg_21__13_ ( .D(n15525), .CK(clk), .RN(rst_n), .Q(
        conv_3[328]) );
  DFFRHQXL conv_3_reg_22__14_ ( .D(n15514), .CK(clk), .RN(rst_n), .Q(
        conv_3[344]) );
  DFFRHQXL conv_3_reg_22__0_ ( .D(n15901), .CK(clk), .RN(rst_n), .Q(
        conv_3[330]) );
  DFFRHQXL conv_3_reg_22__5_ ( .D(n15523), .CK(clk), .RN(rst_n), .Q(
        conv_3[335]) );
  DFFRHQXL conv_3_reg_22__6_ ( .D(n15522), .CK(clk), .RN(rst_n), .Q(
        conv_3[336]) );
  DFFRHQXL conv_3_reg_22__7_ ( .D(n15521), .CK(clk), .RN(rst_n), .Q(
        conv_3[337]) );
  DFFRHQXL conv_3_reg_22__8_ ( .D(n15520), .CK(clk), .RN(rst_n), .Q(
        conv_3[338]) );
  DFFRHQXL conv_3_reg_22__9_ ( .D(n15519), .CK(clk), .RN(rst_n), .Q(
        conv_3[339]) );
  DFFRHQXL conv_3_reg_22__10_ ( .D(n15518), .CK(clk), .RN(rst_n), .Q(
        conv_3[340]) );
  DFFRHQXL conv_3_reg_22__11_ ( .D(n15517), .CK(clk), .RN(rst_n), .Q(
        conv_3[341]) );
  DFFRHQXL conv_3_reg_22__12_ ( .D(n15516), .CK(clk), .RN(rst_n), .Q(
        conv_3[342]) );
  DFFRHQXL conv_3_reg_22__13_ ( .D(n15515), .CK(clk), .RN(rst_n), .Q(
        conv_3[343]) );
  DFFRHQXL conv_3_reg_23__14_ ( .D(n15504), .CK(clk), .RN(rst_n), .Q(
        conv_3[359]) );
  DFFRHQXL conv_3_reg_23__0_ ( .D(n15900), .CK(clk), .RN(rst_n), .Q(
        conv_3[345]) );
  DFFRHQXL conv_3_reg_23__5_ ( .D(n15513), .CK(clk), .RN(rst_n), .Q(
        conv_3[350]) );
  DFFRHQXL conv_3_reg_23__6_ ( .D(n15512), .CK(clk), .RN(rst_n), .Q(
        conv_3[351]) );
  DFFRHQXL conv_3_reg_23__7_ ( .D(n15511), .CK(clk), .RN(rst_n), .Q(
        conv_3[352]) );
  DFFRHQXL conv_3_reg_23__8_ ( .D(n15510), .CK(clk), .RN(rst_n), .Q(
        conv_3[353]) );
  DFFRHQXL conv_3_reg_23__9_ ( .D(n15509), .CK(clk), .RN(rst_n), .Q(
        conv_3[354]) );
  DFFRHQXL conv_3_reg_23__10_ ( .D(n15508), .CK(clk), .RN(rst_n), .Q(
        conv_3[355]) );
  DFFRHQXL conv_3_reg_23__11_ ( .D(n15507), .CK(clk), .RN(rst_n), .Q(
        conv_3[356]) );
  DFFRHQXL conv_3_reg_23__12_ ( .D(n15506), .CK(clk), .RN(rst_n), .Q(
        conv_3[357]) );
  DFFRHQXL conv_3_reg_23__13_ ( .D(n15505), .CK(clk), .RN(rst_n), .Q(
        conv_3[358]) );
  DFFRHQXL conv_3_reg_24__14_ ( .D(n15494), .CK(clk), .RN(rst_n), .Q(
        conv_3[374]) );
  DFFRHQXL conv_3_reg_24__0_ ( .D(n15899), .CK(clk), .RN(rst_n), .Q(
        conv_3[360]) );
  DFFRHQXL conv_3_reg_24__5_ ( .D(n15503), .CK(clk), .RN(rst_n), .Q(
        conv_3[365]) );
  DFFRHQXL conv_3_reg_24__6_ ( .D(n15502), .CK(clk), .RN(rst_n), .Q(
        conv_3[366]) );
  DFFRHQXL conv_3_reg_24__7_ ( .D(n15501), .CK(clk), .RN(rst_n), .Q(
        conv_3[367]) );
  DFFRHQXL conv_3_reg_24__8_ ( .D(n15500), .CK(clk), .RN(rst_n), .Q(
        conv_3[368]) );
  DFFRHQXL conv_3_reg_24__9_ ( .D(n15499), .CK(clk), .RN(rst_n), .Q(
        conv_3[369]) );
  DFFRHQXL conv_3_reg_24__10_ ( .D(n15498), .CK(clk), .RN(rst_n), .Q(
        conv_3[370]) );
  DFFRHQXL conv_3_reg_24__11_ ( .D(n15497), .CK(clk), .RN(rst_n), .Q(
        conv_3[371]) );
  DFFRHQXL conv_3_reg_24__12_ ( .D(n15496), .CK(clk), .RN(rst_n), .Q(
        conv_3[372]) );
  DFFRHQXL conv_3_reg_24__13_ ( .D(n15495), .CK(clk), .RN(rst_n), .Q(
        conv_3[373]) );
  DFFRHQXL conv_3_reg_25__14_ ( .D(n15484), .CK(clk), .RN(rst_n), .Q(
        conv_3[389]) );
  DFFRHQXL conv_3_reg_25__0_ ( .D(n15898), .CK(clk), .RN(rst_n), .Q(
        conv_3[375]) );
  DFFRHQXL conv_3_reg_25__5_ ( .D(n15493), .CK(clk), .RN(rst_n), .Q(
        conv_3[380]) );
  DFFRHQXL conv_3_reg_25__6_ ( .D(n15492), .CK(clk), .RN(rst_n), .Q(
        conv_3[381]) );
  DFFRHQXL conv_3_reg_25__7_ ( .D(n15491), .CK(clk), .RN(rst_n), .Q(
        conv_3[382]) );
  DFFRHQXL conv_3_reg_25__8_ ( .D(n15490), .CK(clk), .RN(rst_n), .Q(
        conv_3[383]) );
  DFFRHQXL conv_3_reg_25__9_ ( .D(n15489), .CK(clk), .RN(rst_n), .Q(
        conv_3[384]) );
  DFFRHQXL conv_3_reg_25__10_ ( .D(n15488), .CK(clk), .RN(rst_n), .Q(
        conv_3[385]) );
  DFFRHQXL conv_3_reg_25__11_ ( .D(n15487), .CK(clk), .RN(rst_n), .Q(
        conv_3[386]) );
  DFFRHQXL conv_3_reg_25__12_ ( .D(n15486), .CK(clk), .RN(rst_n), .Q(
        conv_3[387]) );
  DFFRHQXL conv_3_reg_25__13_ ( .D(n15485), .CK(clk), .RN(rst_n), .Q(
        conv_3[388]) );
  DFFRHQXL conv_3_reg_26__14_ ( .D(n15474), .CK(clk), .RN(rst_n), .Q(
        conv_3[404]) );
  DFFRHQXL conv_3_reg_26__0_ ( .D(n15897), .CK(clk), .RN(rst_n), .Q(
        conv_3[390]) );
  DFFRHQXL conv_3_reg_26__5_ ( .D(n15483), .CK(clk), .RN(rst_n), .Q(
        conv_3[395]) );
  DFFRHQXL conv_3_reg_26__6_ ( .D(n15482), .CK(clk), .RN(rst_n), .Q(
        conv_3[396]) );
  DFFRHQXL conv_3_reg_26__7_ ( .D(n15481), .CK(clk), .RN(rst_n), .Q(
        conv_3[397]) );
  DFFRHQXL conv_3_reg_26__8_ ( .D(n15480), .CK(clk), .RN(rst_n), .Q(
        conv_3[398]) );
  DFFRHQXL conv_3_reg_26__9_ ( .D(n15479), .CK(clk), .RN(rst_n), .Q(
        conv_3[399]) );
  DFFRHQXL conv_3_reg_26__10_ ( .D(n15478), .CK(clk), .RN(rst_n), .Q(
        conv_3[400]) );
  DFFRHQXL conv_3_reg_26__11_ ( .D(n15477), .CK(clk), .RN(rst_n), .Q(
        conv_3[401]) );
  DFFRHQXL conv_3_reg_26__12_ ( .D(n15476), .CK(clk), .RN(rst_n), .Q(
        conv_3[402]) );
  DFFRHQXL conv_3_reg_26__13_ ( .D(n15475), .CK(clk), .RN(rst_n), .Q(
        conv_3[403]) );
  DFFRHQXL conv_3_reg_27__14_ ( .D(n15464), .CK(clk), .RN(rst_n), .Q(
        conv_3[419]) );
  DFFRHQXL conv_3_reg_27__0_ ( .D(n15896), .CK(clk), .RN(rst_n), .Q(
        conv_3[405]) );
  DFFRHQXL conv_3_reg_27__5_ ( .D(n15473), .CK(clk), .RN(rst_n), .Q(
        conv_3[410]) );
  DFFRHQXL conv_3_reg_27__6_ ( .D(n15472), .CK(clk), .RN(rst_n), .Q(
        conv_3[411]) );
  DFFRHQXL conv_3_reg_27__7_ ( .D(n15471), .CK(clk), .RN(rst_n), .Q(
        conv_3[412]) );
  DFFRHQXL conv_3_reg_27__8_ ( .D(n15470), .CK(clk), .RN(rst_n), .Q(
        conv_3[413]) );
  DFFRHQXL conv_3_reg_27__9_ ( .D(n15469), .CK(clk), .RN(rst_n), .Q(
        conv_3[414]) );
  DFFRHQXL conv_3_reg_27__10_ ( .D(n15468), .CK(clk), .RN(rst_n), .Q(
        conv_3[415]) );
  DFFRHQXL conv_3_reg_27__11_ ( .D(n15467), .CK(clk), .RN(rst_n), .Q(
        conv_3[416]) );
  DFFRHQXL conv_3_reg_27__12_ ( .D(n15466), .CK(clk), .RN(rst_n), .Q(
        conv_3[417]) );
  DFFRHQXL conv_3_reg_27__13_ ( .D(n15465), .CK(clk), .RN(rst_n), .Q(
        conv_3[418]) );
  DFFRHQXL conv_3_reg_28__14_ ( .D(n15454), .CK(clk), .RN(rst_n), .Q(
        conv_3[434]) );
  DFFRHQXL conv_3_reg_28__0_ ( .D(n15895), .CK(clk), .RN(rst_n), .Q(
        conv_3[420]) );
  DFFRHQXL conv_3_reg_28__5_ ( .D(n15463), .CK(clk), .RN(rst_n), .Q(
        conv_3[425]) );
  DFFRHQXL conv_3_reg_28__6_ ( .D(n15462), .CK(clk), .RN(rst_n), .Q(
        conv_3[426]) );
  DFFRHQXL conv_3_reg_28__7_ ( .D(n15461), .CK(clk), .RN(rst_n), .Q(
        conv_3[427]) );
  DFFRHQXL conv_3_reg_28__8_ ( .D(n15460), .CK(clk), .RN(rst_n), .Q(
        conv_3[428]) );
  DFFRHQXL conv_3_reg_28__9_ ( .D(n15459), .CK(clk), .RN(rst_n), .Q(
        conv_3[429]) );
  DFFRHQXL conv_3_reg_28__10_ ( .D(n15458), .CK(clk), .RN(rst_n), .Q(
        conv_3[430]) );
  DFFRHQXL conv_3_reg_28__11_ ( .D(n15457), .CK(clk), .RN(rst_n), .Q(
        conv_3[431]) );
  DFFRHQXL conv_3_reg_28__12_ ( .D(n15456), .CK(clk), .RN(rst_n), .Q(
        conv_3[432]) );
  DFFRHQXL conv_3_reg_28__13_ ( .D(n15455), .CK(clk), .RN(rst_n), .Q(
        conv_3[433]) );
  DFFRHQXL conv_3_reg_29__14_ ( .D(n15444), .CK(clk), .RN(rst_n), .Q(
        conv_3[449]) );
  DFFRHQXL conv_3_reg_29__0_ ( .D(n15894), .CK(clk), .RN(rst_n), .Q(
        conv_3[435]) );
  DFFRHQXL conv_3_reg_29__5_ ( .D(n15453), .CK(clk), .RN(rst_n), .Q(
        conv_3[440]) );
  DFFRHQXL conv_3_reg_29__6_ ( .D(n15452), .CK(clk), .RN(rst_n), .Q(
        conv_3[441]) );
  DFFRHQXL conv_3_reg_29__7_ ( .D(n15451), .CK(clk), .RN(rst_n), .Q(
        conv_3[442]) );
  DFFRHQXL conv_3_reg_29__8_ ( .D(n15450), .CK(clk), .RN(rst_n), .Q(
        conv_3[443]) );
  DFFRHQXL conv_3_reg_29__9_ ( .D(n15449), .CK(clk), .RN(rst_n), .Q(
        conv_3[444]) );
  DFFRHQXL conv_3_reg_29__10_ ( .D(n15448), .CK(clk), .RN(rst_n), .Q(
        conv_3[445]) );
  DFFRHQXL conv_3_reg_29__11_ ( .D(n15447), .CK(clk), .RN(rst_n), .Q(
        conv_3[446]) );
  DFFRHQXL conv_3_reg_29__12_ ( .D(n15446), .CK(clk), .RN(rst_n), .Q(
        conv_3[447]) );
  DFFRHQXL conv_3_reg_29__13_ ( .D(n15445), .CK(clk), .RN(rst_n), .Q(
        conv_3[448]) );
  DFFRHQXL conv_3_reg_30__14_ ( .D(n15434), .CK(clk), .RN(rst_n), .Q(
        conv_3[464]) );
  DFFRHQXL conv_3_reg_30__0_ ( .D(n15893), .CK(clk), .RN(rst_n), .Q(
        conv_3[450]) );
  DFFRHQXL conv_3_reg_30__5_ ( .D(n15443), .CK(clk), .RN(rst_n), .Q(
        conv_3[455]) );
  DFFRHQXL conv_3_reg_30__6_ ( .D(n15442), .CK(clk), .RN(rst_n), .Q(
        conv_3[456]) );
  DFFRHQXL conv_3_reg_30__7_ ( .D(n15441), .CK(clk), .RN(rst_n), .Q(
        conv_3[457]) );
  DFFRHQXL conv_3_reg_30__8_ ( .D(n15440), .CK(clk), .RN(rst_n), .Q(
        conv_3[458]) );
  DFFRHQXL conv_3_reg_30__9_ ( .D(n15439), .CK(clk), .RN(rst_n), .Q(
        conv_3[459]) );
  DFFRHQXL conv_3_reg_30__10_ ( .D(n15438), .CK(clk), .RN(rst_n), .Q(
        conv_3[460]) );
  DFFRHQXL conv_3_reg_30__11_ ( .D(n15437), .CK(clk), .RN(rst_n), .Q(
        conv_3[461]) );
  DFFRHQXL conv_3_reg_30__12_ ( .D(n15436), .CK(clk), .RN(rst_n), .Q(
        conv_3[462]) );
  DFFRHQXL conv_3_reg_30__13_ ( .D(n15435), .CK(clk), .RN(rst_n), .Q(
        conv_3[463]) );
  DFFRHQXL conv_3_reg_31__14_ ( .D(n15424), .CK(clk), .RN(rst_n), .Q(
        conv_3[479]) );
  DFFRHQXL conv_3_reg_31__0_ ( .D(n15892), .CK(clk), .RN(rst_n), .Q(
        conv_3[465]) );
  DFFRHQXL conv_3_reg_31__5_ ( .D(n15433), .CK(clk), .RN(rst_n), .Q(
        conv_3[470]) );
  DFFRHQXL conv_3_reg_31__6_ ( .D(n15432), .CK(clk), .RN(rst_n), .Q(
        conv_3[471]) );
  DFFRHQXL conv_3_reg_31__7_ ( .D(n15431), .CK(clk), .RN(rst_n), .Q(
        conv_3[472]) );
  DFFRHQXL conv_3_reg_31__8_ ( .D(n15430), .CK(clk), .RN(rst_n), .Q(
        conv_3[473]) );
  DFFRHQXL conv_3_reg_31__9_ ( .D(n15429), .CK(clk), .RN(rst_n), .Q(
        conv_3[474]) );
  DFFRHQXL conv_3_reg_31__10_ ( .D(n15428), .CK(clk), .RN(rst_n), .Q(
        conv_3[475]) );
  DFFRHQXL conv_3_reg_31__11_ ( .D(n15427), .CK(clk), .RN(rst_n), .Q(
        conv_3[476]) );
  DFFRHQXL conv_3_reg_31__12_ ( .D(n15426), .CK(clk), .RN(rst_n), .Q(
        conv_3[477]) );
  DFFRHQXL conv_3_reg_31__13_ ( .D(n15425), .CK(clk), .RN(rst_n), .Q(
        conv_3[478]) );
  DFFRHQXL conv_3_reg_32__14_ ( .D(n15414), .CK(clk), .RN(rst_n), .Q(
        conv_3[494]) );
  DFFRHQXL conv_3_reg_32__0_ ( .D(n15891), .CK(clk), .RN(rst_n), .Q(
        conv_3[480]) );
  DFFRHQXL conv_3_reg_32__5_ ( .D(n15423), .CK(clk), .RN(rst_n), .Q(
        conv_3[485]) );
  DFFRHQXL conv_3_reg_32__6_ ( .D(n15422), .CK(clk), .RN(rst_n), .Q(
        conv_3[486]) );
  DFFRHQXL conv_3_reg_32__7_ ( .D(n15421), .CK(clk), .RN(rst_n), .Q(
        conv_3[487]) );
  DFFRHQXL conv_3_reg_32__8_ ( .D(n15420), .CK(clk), .RN(rst_n), .Q(
        conv_3[488]) );
  DFFRHQXL conv_3_reg_32__9_ ( .D(n15419), .CK(clk), .RN(rst_n), .Q(
        conv_3[489]) );
  DFFRHQXL conv_3_reg_32__10_ ( .D(n15418), .CK(clk), .RN(rst_n), .Q(
        conv_3[490]) );
  DFFRHQXL conv_3_reg_32__11_ ( .D(n15417), .CK(clk), .RN(rst_n), .Q(
        conv_3[491]) );
  DFFRHQXL conv_3_reg_32__12_ ( .D(n15416), .CK(clk), .RN(rst_n), .Q(
        conv_3[492]) );
  DFFRHQXL conv_3_reg_32__13_ ( .D(n15415), .CK(clk), .RN(rst_n), .Q(
        conv_3[493]) );
  DFFRHQXL conv_3_reg_33__14_ ( .D(n15404), .CK(clk), .RN(rst_n), .Q(
        conv_3[509]) );
  DFFRHQXL conv_3_reg_33__0_ ( .D(n15890), .CK(clk), .RN(rst_n), .Q(
        conv_3[495]) );
  DFFRHQXL conv_3_reg_33__5_ ( .D(n15413), .CK(clk), .RN(rst_n), .Q(
        conv_3[500]) );
  DFFRHQXL conv_3_reg_33__6_ ( .D(n15412), .CK(clk), .RN(rst_n), .Q(
        conv_3[501]) );
  DFFRHQXL conv_3_reg_33__7_ ( .D(n15411), .CK(clk), .RN(rst_n), .Q(
        conv_3[502]) );
  DFFRHQXL conv_3_reg_33__8_ ( .D(n15410), .CK(clk), .RN(rst_n), .Q(
        conv_3[503]) );
  DFFRHQXL conv_3_reg_33__9_ ( .D(n15409), .CK(clk), .RN(rst_n), .Q(
        conv_3[504]) );
  DFFRHQXL conv_3_reg_33__10_ ( .D(n15408), .CK(clk), .RN(rst_n), .Q(
        conv_3[505]) );
  DFFRHQXL conv_3_reg_33__11_ ( .D(n15407), .CK(clk), .RN(rst_n), .Q(
        conv_3[506]) );
  DFFRHQXL conv_3_reg_33__12_ ( .D(n15406), .CK(clk), .RN(rst_n), .Q(
        conv_3[507]) );
  DFFRHQXL conv_3_reg_33__13_ ( .D(n15405), .CK(clk), .RN(rst_n), .Q(
        conv_3[508]) );
  DFFRHQXL conv_3_reg_34__14_ ( .D(n15394), .CK(clk), .RN(rst_n), .Q(
        conv_3[524]) );
  DFFRHQXL conv_3_reg_34__0_ ( .D(n15889), .CK(clk), .RN(rst_n), .Q(
        conv_3[510]) );
  DFFRHQXL conv_3_reg_34__5_ ( .D(n15403), .CK(clk), .RN(rst_n), .Q(
        conv_3[515]) );
  DFFRHQXL conv_3_reg_34__6_ ( .D(n15402), .CK(clk), .RN(rst_n), .Q(
        conv_3[516]) );
  DFFRHQXL conv_3_reg_34__7_ ( .D(n15401), .CK(clk), .RN(rst_n), .Q(
        conv_3[517]) );
  DFFRHQXL conv_3_reg_34__8_ ( .D(n15400), .CK(clk), .RN(rst_n), .Q(
        conv_3[518]) );
  DFFRHQXL conv_3_reg_34__9_ ( .D(n15399), .CK(clk), .RN(rst_n), .Q(
        conv_3[519]) );
  DFFRHQXL conv_3_reg_34__10_ ( .D(n15398), .CK(clk), .RN(rst_n), .Q(
        conv_3[520]) );
  DFFRHQXL conv_3_reg_34__11_ ( .D(n15397), .CK(clk), .RN(rst_n), .Q(
        conv_3[521]) );
  DFFRHQXL conv_3_reg_34__12_ ( .D(n15396), .CK(clk), .RN(rst_n), .Q(
        conv_3[522]) );
  DFFRHQXL conv_3_reg_34__13_ ( .D(n15395), .CK(clk), .RN(rst_n), .Q(
        conv_3[523]) );
  DFFRHQXL conv_3_reg_35__14_ ( .D(n15384), .CK(clk), .RN(rst_n), .Q(
        conv_3[539]) );
  DFFRHQXL conv_3_reg_35__0_ ( .D(n15888), .CK(clk), .RN(rst_n), .Q(
        conv_3[525]) );
  DFFRHQXL pool_reg_24__0_ ( .D(N29336), .CK(clk), .RN(rst_n), .Q(pool[120])
         );
  DFFRHQXL pool_reg_26__0_ ( .D(N29346), .CK(clk), .RN(rst_n), .Q(pool[130])
         );
  DFFRHQXL pool_reg_21__0_ ( .D(N29321), .CK(clk), .RN(rst_n), .Q(pool[105])
         );
  DFFRHQXL pool_reg_20__0_ ( .D(N29316), .CK(clk), .RN(rst_n), .Q(pool[100])
         );
  DFFRHQXL pool_reg_23__0_ ( .D(N29331), .CK(clk), .RN(rst_n), .Q(pool[115])
         );
  DFFRHQXL pool_reg_18__0_ ( .D(N29306), .CK(clk), .RN(rst_n), .Q(pool[90]) );
  DFFRHQXL pool_reg_19__0_ ( .D(N29311), .CK(clk), .RN(rst_n), .Q(pool[95]) );
  DFFRHQXL pool_reg_25__0_ ( .D(N29341), .CK(clk), .RN(rst_n), .Q(pool[125])
         );
  DFFRHQXL pool_reg_22__0_ ( .D(N29326), .CK(clk), .RN(rst_n), .Q(pool[110])
         );
  DFFRHQXL conv_3_reg_35__5_ ( .D(n15393), .CK(clk), .RN(rst_n), .Q(
        conv_3[530]) );
  DFFRHQXL conv_3_reg_35__6_ ( .D(n15392), .CK(clk), .RN(rst_n), .Q(
        conv_3[531]) );
  DFFRHQXL conv_3_reg_35__7_ ( .D(n15391), .CK(clk), .RN(rst_n), .Q(
        conv_3[532]) );
  DFFRHQXL conv_3_reg_35__8_ ( .D(n15390), .CK(clk), .RN(rst_n), .Q(
        conv_3[533]) );
  DFFRHQXL conv_3_reg_35__9_ ( .D(n15389), .CK(clk), .RN(rst_n), .Q(
        conv_3[534]) );
  DFFRHQXL conv_3_reg_35__10_ ( .D(n15388), .CK(clk), .RN(rst_n), .Q(
        conv_3[535]) );
  DFFRHQXL conv_3_reg_35__11_ ( .D(n15387), .CK(clk), .RN(rst_n), .Q(
        conv_3[536]) );
  DFFRHQXL conv_3_reg_35__12_ ( .D(n15386), .CK(clk), .RN(rst_n), .Q(
        conv_3[537]) );
  DFFRHQXL conv_3_reg_35__13_ ( .D(n15385), .CK(clk), .RN(rst_n), .Q(
        conv_3[538]) );
  DFFRHQXL filter_2_bias_reg_5_ ( .D(n14731), .CK(clk), .RN(rst_n), .Q(
        filter_2_bias[5]) );
  DFFRHQXL conv_2_reg_0__14_ ( .D(n15194), .CK(clk), .RN(rst_n), .Q(conv_2[14]) );
  DFFRHQXL conv_2_reg_0__0_ ( .D(n15383), .CK(clk), .RN(rst_n), .Q(conv_2[0])
         );
  DFFRHQXL conv_2_reg_0__5_ ( .D(n15203), .CK(clk), .RN(rst_n), .Q(conv_2[5])
         );
  DFFRHQXL conv_2_reg_0__6_ ( .D(n15202), .CK(clk), .RN(rst_n), .Q(conv_2[6])
         );
  DFFRHQXL conv_2_reg_0__7_ ( .D(n15201), .CK(clk), .RN(rst_n), .Q(conv_2[7])
         );
  DFFRHQXL conv_2_reg_0__8_ ( .D(n15200), .CK(clk), .RN(rst_n), .Q(conv_2[8])
         );
  DFFRHQXL conv_2_reg_0__9_ ( .D(n15199), .CK(clk), .RN(rst_n), .Q(conv_2[9])
         );
  DFFRHQXL conv_2_reg_0__10_ ( .D(n15198), .CK(clk), .RN(rst_n), .Q(conv_2[10]) );
  DFFRHQXL conv_2_reg_0__11_ ( .D(n15197), .CK(clk), .RN(rst_n), .Q(conv_2[11]) );
  DFFRHQXL conv_2_reg_0__12_ ( .D(n15196), .CK(clk), .RN(rst_n), .Q(conv_2[12]) );
  DFFRHQXL conv_2_reg_0__13_ ( .D(n15195), .CK(clk), .RN(rst_n), .Q(conv_2[13]) );
  DFFRHQXL conv_2_reg_1__14_ ( .D(n15184), .CK(clk), .RN(rst_n), .Q(conv_2[29]) );
  DFFRHQXL conv_2_reg_1__0_ ( .D(n15382), .CK(clk), .RN(rst_n), .Q(conv_2[15])
         );
  DFFRHQXL conv_2_reg_1__5_ ( .D(n15193), .CK(clk), .RN(rst_n), .Q(conv_2[20])
         );
  DFFRHQXL conv_2_reg_1__6_ ( .D(n15192), .CK(clk), .RN(rst_n), .Q(conv_2[21])
         );
  DFFRHQXL conv_2_reg_1__7_ ( .D(n15191), .CK(clk), .RN(rst_n), .Q(conv_2[22])
         );
  DFFRHQXL conv_2_reg_1__8_ ( .D(n15190), .CK(clk), .RN(rst_n), .Q(conv_2[23])
         );
  DFFRHQXL conv_2_reg_1__9_ ( .D(n15189), .CK(clk), .RN(rst_n), .Q(conv_2[24])
         );
  DFFRHQXL conv_2_reg_1__10_ ( .D(n15188), .CK(clk), .RN(rst_n), .Q(conv_2[25]) );
  DFFRHQXL conv_2_reg_1__11_ ( .D(n15187), .CK(clk), .RN(rst_n), .Q(conv_2[26]) );
  DFFRHQXL conv_2_reg_1__12_ ( .D(n15186), .CK(clk), .RN(rst_n), .Q(conv_2[27]) );
  DFFRHQXL conv_2_reg_1__13_ ( .D(n15185), .CK(clk), .RN(rst_n), .Q(conv_2[28]) );
  DFFRHQXL conv_2_reg_2__14_ ( .D(n15174), .CK(clk), .RN(rst_n), .Q(conv_2[44]) );
  DFFRHQXL conv_2_reg_2__0_ ( .D(n15381), .CK(clk), .RN(rst_n), .Q(conv_2[30])
         );
  DFFRHQXL conv_2_reg_2__5_ ( .D(n15183), .CK(clk), .RN(rst_n), .Q(conv_2[35])
         );
  DFFRHQXL conv_2_reg_2__6_ ( .D(n15182), .CK(clk), .RN(rst_n), .Q(conv_2[36])
         );
  DFFRHQXL conv_2_reg_2__7_ ( .D(n15181), .CK(clk), .RN(rst_n), .Q(conv_2[37])
         );
  DFFRHQXL conv_2_reg_2__8_ ( .D(n15180), .CK(clk), .RN(rst_n), .Q(conv_2[38])
         );
  DFFRHQXL conv_2_reg_2__9_ ( .D(n15179), .CK(clk), .RN(rst_n), .Q(conv_2[39])
         );
  DFFRHQXL conv_2_reg_2__10_ ( .D(n15178), .CK(clk), .RN(rst_n), .Q(conv_2[40]) );
  DFFRHQXL conv_2_reg_2__11_ ( .D(n15177), .CK(clk), .RN(rst_n), .Q(conv_2[41]) );
  DFFRHQXL conv_2_reg_2__12_ ( .D(n15176), .CK(clk), .RN(rst_n), .Q(conv_2[42]) );
  DFFRHQXL conv_2_reg_2__13_ ( .D(n15175), .CK(clk), .RN(rst_n), .Q(conv_2[43]) );
  DFFRHQXL conv_2_reg_3__14_ ( .D(n15164), .CK(clk), .RN(rst_n), .Q(conv_2[59]) );
  DFFRHQXL conv_2_reg_3__0_ ( .D(n15380), .CK(clk), .RN(rst_n), .Q(conv_2[45])
         );
  DFFRHQXL conv_2_reg_3__5_ ( .D(n15173), .CK(clk), .RN(rst_n), .Q(conv_2[50])
         );
  DFFRHQXL conv_2_reg_3__6_ ( .D(n15172), .CK(clk), .RN(rst_n), .Q(conv_2[51])
         );
  DFFRHQXL conv_2_reg_3__7_ ( .D(n15171), .CK(clk), .RN(rst_n), .Q(conv_2[52])
         );
  DFFRHQXL conv_2_reg_3__8_ ( .D(n15170), .CK(clk), .RN(rst_n), .Q(conv_2[53])
         );
  DFFRHQXL conv_2_reg_3__9_ ( .D(n15169), .CK(clk), .RN(rst_n), .Q(conv_2[54])
         );
  DFFRHQXL conv_2_reg_3__10_ ( .D(n15168), .CK(clk), .RN(rst_n), .Q(conv_2[55]) );
  DFFRHQXL conv_2_reg_3__11_ ( .D(n15167), .CK(clk), .RN(rst_n), .Q(conv_2[56]) );
  DFFRHQXL conv_2_reg_3__12_ ( .D(n15166), .CK(clk), .RN(rst_n), .Q(conv_2[57]) );
  DFFRHQXL conv_2_reg_3__13_ ( .D(n15165), .CK(clk), .RN(rst_n), .Q(conv_2[58]) );
  DFFRHQXL conv_2_reg_4__14_ ( .D(n15154), .CK(clk), .RN(rst_n), .Q(conv_2[74]) );
  DFFRHQXL conv_2_reg_4__0_ ( .D(n15379), .CK(clk), .RN(rst_n), .Q(conv_2[60])
         );
  DFFRHQXL conv_2_reg_4__5_ ( .D(n15163), .CK(clk), .RN(rst_n), .Q(conv_2[65])
         );
  DFFRHQXL conv_2_reg_4__6_ ( .D(n15162), .CK(clk), .RN(rst_n), .Q(conv_2[66])
         );
  DFFRHQXL conv_2_reg_4__7_ ( .D(n15161), .CK(clk), .RN(rst_n), .Q(conv_2[67])
         );
  DFFRHQXL conv_2_reg_4__8_ ( .D(n15160), .CK(clk), .RN(rst_n), .Q(conv_2[68])
         );
  DFFRHQXL conv_2_reg_4__9_ ( .D(n15159), .CK(clk), .RN(rst_n), .Q(conv_2[69])
         );
  DFFRHQXL conv_2_reg_4__10_ ( .D(n15158), .CK(clk), .RN(rst_n), .Q(conv_2[70]) );
  DFFRHQXL conv_2_reg_4__11_ ( .D(n15157), .CK(clk), .RN(rst_n), .Q(conv_2[71]) );
  DFFRHQXL conv_2_reg_4__12_ ( .D(n15156), .CK(clk), .RN(rst_n), .Q(conv_2[72]) );
  DFFRHQXL conv_2_reg_4__13_ ( .D(n15155), .CK(clk), .RN(rst_n), .Q(conv_2[73]) );
  DFFRHQXL conv_2_reg_5__14_ ( .D(n15144), .CK(clk), .RN(rst_n), .Q(conv_2[89]) );
  DFFRHQXL conv_2_reg_5__0_ ( .D(n15378), .CK(clk), .RN(rst_n), .Q(conv_2[75])
         );
  DFFRHQXL conv_2_reg_5__5_ ( .D(n15153), .CK(clk), .RN(rst_n), .Q(conv_2[80])
         );
  DFFRHQXL conv_2_reg_5__6_ ( .D(n15152), .CK(clk), .RN(rst_n), .Q(conv_2[81])
         );
  DFFRHQXL conv_2_reg_5__7_ ( .D(n15151), .CK(clk), .RN(rst_n), .Q(conv_2[82])
         );
  DFFRHQXL conv_2_reg_5__8_ ( .D(n15150), .CK(clk), .RN(rst_n), .Q(conv_2[83])
         );
  DFFRHQXL conv_2_reg_5__9_ ( .D(n15149), .CK(clk), .RN(rst_n), .Q(conv_2[84])
         );
  DFFRHQXL conv_2_reg_5__10_ ( .D(n15148), .CK(clk), .RN(rst_n), .Q(conv_2[85]) );
  DFFRHQXL conv_2_reg_5__11_ ( .D(n15147), .CK(clk), .RN(rst_n), .Q(conv_2[86]) );
  DFFRHQXL conv_2_reg_5__12_ ( .D(n15146), .CK(clk), .RN(rst_n), .Q(conv_2[87]) );
  DFFRHQXL conv_2_reg_5__13_ ( .D(n15145), .CK(clk), .RN(rst_n), .Q(conv_2[88]) );
  DFFRHQXL conv_2_reg_6__14_ ( .D(n15134), .CK(clk), .RN(rst_n), .Q(
        conv_2[104]) );
  DFFRHQXL conv_2_reg_6__0_ ( .D(n15377), .CK(clk), .RN(rst_n), .Q(conv_2[90])
         );
  DFFRHQXL conv_2_reg_6__5_ ( .D(n15143), .CK(clk), .RN(rst_n), .Q(conv_2[95])
         );
  DFFRHQXL conv_2_reg_6__6_ ( .D(n15142), .CK(clk), .RN(rst_n), .Q(conv_2[96])
         );
  DFFRHQXL conv_2_reg_6__7_ ( .D(n15141), .CK(clk), .RN(rst_n), .Q(conv_2[97])
         );
  DFFRHQXL conv_2_reg_6__8_ ( .D(n15140), .CK(clk), .RN(rst_n), .Q(conv_2[98])
         );
  DFFRHQXL conv_2_reg_6__9_ ( .D(n15139), .CK(clk), .RN(rst_n), .Q(conv_2[99])
         );
  DFFRHQXL conv_2_reg_6__10_ ( .D(n15138), .CK(clk), .RN(rst_n), .Q(
        conv_2[100]) );
  DFFRHQXL conv_2_reg_6__11_ ( .D(n15137), .CK(clk), .RN(rst_n), .Q(
        conv_2[101]) );
  DFFRHQXL conv_2_reg_6__12_ ( .D(n15136), .CK(clk), .RN(rst_n), .Q(
        conv_2[102]) );
  DFFRHQXL conv_2_reg_6__13_ ( .D(n15135), .CK(clk), .RN(rst_n), .Q(
        conv_2[103]) );
  DFFRHQXL conv_2_reg_7__14_ ( .D(n15124), .CK(clk), .RN(rst_n), .Q(
        conv_2[119]) );
  DFFRHQXL conv_2_reg_7__0_ ( .D(n15376), .CK(clk), .RN(rst_n), .Q(conv_2[105]) );
  DFFRHQXL conv_2_reg_7__5_ ( .D(n15133), .CK(clk), .RN(rst_n), .Q(conv_2[110]) );
  DFFRHQXL conv_2_reg_7__6_ ( .D(n15132), .CK(clk), .RN(rst_n), .Q(conv_2[111]) );
  DFFRHQXL conv_2_reg_7__7_ ( .D(n15131), .CK(clk), .RN(rst_n), .Q(conv_2[112]) );
  DFFRHQXL conv_2_reg_7__8_ ( .D(n15130), .CK(clk), .RN(rst_n), .Q(conv_2[113]) );
  DFFRHQXL conv_2_reg_7__9_ ( .D(n15129), .CK(clk), .RN(rst_n), .Q(conv_2[114]) );
  DFFRHQXL conv_2_reg_7__10_ ( .D(n15128), .CK(clk), .RN(rst_n), .Q(
        conv_2[115]) );
  DFFRHQXL conv_2_reg_7__11_ ( .D(n15127), .CK(clk), .RN(rst_n), .Q(
        conv_2[116]) );
  DFFRHQXL conv_2_reg_7__12_ ( .D(n15126), .CK(clk), .RN(rst_n), .Q(
        conv_2[117]) );
  DFFRHQXL conv_2_reg_7__13_ ( .D(n15125), .CK(clk), .RN(rst_n), .Q(
        conv_2[118]) );
  DFFRHQXL conv_2_reg_8__14_ ( .D(n15114), .CK(clk), .RN(rst_n), .Q(
        conv_2[134]) );
  DFFRHQXL conv_2_reg_8__0_ ( .D(n15375), .CK(clk), .RN(rst_n), .Q(conv_2[120]) );
  DFFRHQXL conv_2_reg_8__5_ ( .D(n15123), .CK(clk), .RN(rst_n), .Q(conv_2[125]) );
  DFFRHQXL conv_2_reg_8__6_ ( .D(n15122), .CK(clk), .RN(rst_n), .Q(conv_2[126]) );
  DFFRHQXL conv_2_reg_8__7_ ( .D(n15121), .CK(clk), .RN(rst_n), .Q(conv_2[127]) );
  DFFRHQXL conv_2_reg_8__8_ ( .D(n15120), .CK(clk), .RN(rst_n), .Q(conv_2[128]) );
  DFFRHQXL conv_2_reg_8__9_ ( .D(n15119), .CK(clk), .RN(rst_n), .Q(conv_2[129]) );
  DFFRHQXL conv_2_reg_8__10_ ( .D(n15118), .CK(clk), .RN(rst_n), .Q(
        conv_2[130]) );
  DFFRHQXL conv_2_reg_8__11_ ( .D(n15117), .CK(clk), .RN(rst_n), .Q(
        conv_2[131]) );
  DFFRHQXL conv_2_reg_8__12_ ( .D(n15116), .CK(clk), .RN(rst_n), .Q(
        conv_2[132]) );
  DFFRHQXL conv_2_reg_8__13_ ( .D(n15115), .CK(clk), .RN(rst_n), .Q(
        conv_2[133]) );
  DFFRHQXL conv_2_reg_9__14_ ( .D(n15104), .CK(clk), .RN(rst_n), .Q(
        conv_2[149]) );
  DFFRHQXL conv_2_reg_9__0_ ( .D(n15374), .CK(clk), .RN(rst_n), .Q(conv_2[135]) );
  DFFRHQXL conv_2_reg_9__5_ ( .D(n15113), .CK(clk), .RN(rst_n), .Q(conv_2[140]) );
  DFFRHQXL conv_2_reg_9__6_ ( .D(n15112), .CK(clk), .RN(rst_n), .Q(conv_2[141]) );
  DFFRHQXL conv_2_reg_9__7_ ( .D(n15111), .CK(clk), .RN(rst_n), .Q(conv_2[142]) );
  DFFRHQXL conv_2_reg_9__8_ ( .D(n15110), .CK(clk), .RN(rst_n), .Q(conv_2[143]) );
  DFFRHQXL conv_2_reg_9__9_ ( .D(n15109), .CK(clk), .RN(rst_n), .Q(conv_2[144]) );
  DFFRHQXL conv_2_reg_9__10_ ( .D(n15108), .CK(clk), .RN(rst_n), .Q(
        conv_2[145]) );
  DFFRHQXL conv_2_reg_9__11_ ( .D(n15107), .CK(clk), .RN(rst_n), .Q(
        conv_2[146]) );
  DFFRHQXL conv_2_reg_9__12_ ( .D(n15106), .CK(clk), .RN(rst_n), .Q(
        conv_2[147]) );
  DFFRHQXL conv_2_reg_9__13_ ( .D(n15105), .CK(clk), .RN(rst_n), .Q(
        conv_2[148]) );
  DFFRHQXL conv_2_reg_10__14_ ( .D(n15094), .CK(clk), .RN(rst_n), .Q(
        conv_2[164]) );
  DFFRHQXL conv_2_reg_10__0_ ( .D(n15373), .CK(clk), .RN(rst_n), .Q(
        conv_2[150]) );
  DFFRHQXL conv_2_reg_10__5_ ( .D(n15103), .CK(clk), .RN(rst_n), .Q(
        conv_2[155]) );
  DFFRHQXL conv_2_reg_10__6_ ( .D(n15102), .CK(clk), .RN(rst_n), .Q(
        conv_2[156]) );
  DFFRHQXL conv_2_reg_10__7_ ( .D(n15101), .CK(clk), .RN(rst_n), .Q(
        conv_2[157]) );
  DFFRHQXL conv_2_reg_10__8_ ( .D(n15100), .CK(clk), .RN(rst_n), .Q(
        conv_2[158]) );
  DFFRHQXL conv_2_reg_10__9_ ( .D(n15099), .CK(clk), .RN(rst_n), .Q(
        conv_2[159]) );
  DFFRHQXL conv_2_reg_10__10_ ( .D(n15098), .CK(clk), .RN(rst_n), .Q(
        conv_2[160]) );
  DFFRHQXL conv_2_reg_10__11_ ( .D(n15097), .CK(clk), .RN(rst_n), .Q(
        conv_2[161]) );
  DFFRHQXL conv_2_reg_10__12_ ( .D(n15096), .CK(clk), .RN(rst_n), .Q(
        conv_2[162]) );
  DFFRHQXL conv_2_reg_10__13_ ( .D(n15095), .CK(clk), .RN(rst_n), .Q(
        conv_2[163]) );
  DFFRHQXL conv_2_reg_11__14_ ( .D(n15084), .CK(clk), .RN(rst_n), .Q(
        conv_2[179]) );
  DFFRHQXL conv_2_reg_11__0_ ( .D(n15372), .CK(clk), .RN(rst_n), .Q(
        conv_2[165]) );
  DFFRHQXL conv_2_reg_11__5_ ( .D(n15093), .CK(clk), .RN(rst_n), .Q(
        conv_2[170]) );
  DFFRHQXL conv_2_reg_11__6_ ( .D(n15092), .CK(clk), .RN(rst_n), .Q(
        conv_2[171]) );
  DFFRHQXL conv_2_reg_11__7_ ( .D(n15091), .CK(clk), .RN(rst_n), .Q(
        conv_2[172]) );
  DFFRHQXL conv_2_reg_11__8_ ( .D(n15090), .CK(clk), .RN(rst_n), .Q(
        conv_2[173]) );
  DFFRHQXL conv_2_reg_11__9_ ( .D(n15089), .CK(clk), .RN(rst_n), .Q(
        conv_2[174]) );
  DFFRHQXL conv_2_reg_11__10_ ( .D(n15088), .CK(clk), .RN(rst_n), .Q(
        conv_2[175]) );
  DFFRHQXL conv_2_reg_11__11_ ( .D(n15087), .CK(clk), .RN(rst_n), .Q(
        conv_2[176]) );
  DFFRHQXL conv_2_reg_11__12_ ( .D(n15086), .CK(clk), .RN(rst_n), .Q(
        conv_2[177]) );
  DFFRHQXL conv_2_reg_11__13_ ( .D(n15085), .CK(clk), .RN(rst_n), .Q(
        conv_2[178]) );
  DFFRHQXL conv_2_reg_12__14_ ( .D(n15074), .CK(clk), .RN(rst_n), .Q(
        conv_2[194]) );
  DFFRHQXL conv_2_reg_12__0_ ( .D(n15371), .CK(clk), .RN(rst_n), .Q(
        conv_2[180]) );
  DFFRHQXL conv_2_reg_12__5_ ( .D(n15083), .CK(clk), .RN(rst_n), .Q(
        conv_2[185]) );
  DFFRHQXL conv_2_reg_12__6_ ( .D(n15082), .CK(clk), .RN(rst_n), .Q(
        conv_2[186]) );
  DFFRHQXL conv_2_reg_12__7_ ( .D(n15081), .CK(clk), .RN(rst_n), .Q(
        conv_2[187]) );
  DFFRHQXL conv_2_reg_12__8_ ( .D(n15080), .CK(clk), .RN(rst_n), .Q(
        conv_2[188]) );
  DFFRHQXL conv_2_reg_12__9_ ( .D(n15079), .CK(clk), .RN(rst_n), .Q(
        conv_2[189]) );
  DFFRHQXL conv_2_reg_12__10_ ( .D(n15078), .CK(clk), .RN(rst_n), .Q(
        conv_2[190]) );
  DFFRHQXL conv_2_reg_12__11_ ( .D(n15077), .CK(clk), .RN(rst_n), .Q(
        conv_2[191]) );
  DFFRHQXL conv_2_reg_12__12_ ( .D(n15076), .CK(clk), .RN(rst_n), .Q(
        conv_2[192]) );
  DFFRHQXL conv_2_reg_12__13_ ( .D(n15075), .CK(clk), .RN(rst_n), .Q(
        conv_2[193]) );
  DFFRHQXL conv_2_reg_13__14_ ( .D(n15064), .CK(clk), .RN(rst_n), .Q(
        conv_2[209]) );
  DFFRHQXL conv_2_reg_13__0_ ( .D(n15370), .CK(clk), .RN(rst_n), .Q(
        conv_2[195]) );
  DFFRHQXL conv_2_reg_13__5_ ( .D(n15073), .CK(clk), .RN(rst_n), .Q(
        conv_2[200]) );
  DFFRHQXL conv_2_reg_13__6_ ( .D(n15072), .CK(clk), .RN(rst_n), .Q(
        conv_2[201]) );
  DFFRHQXL conv_2_reg_13__7_ ( .D(n15071), .CK(clk), .RN(rst_n), .Q(
        conv_2[202]) );
  DFFRHQXL conv_2_reg_13__8_ ( .D(n15070), .CK(clk), .RN(rst_n), .Q(
        conv_2[203]) );
  DFFRHQXL conv_2_reg_13__9_ ( .D(n15069), .CK(clk), .RN(rst_n), .Q(
        conv_2[204]) );
  DFFRHQXL conv_2_reg_13__10_ ( .D(n15068), .CK(clk), .RN(rst_n), .Q(
        conv_2[205]) );
  DFFRHQXL conv_2_reg_13__11_ ( .D(n15067), .CK(clk), .RN(rst_n), .Q(
        conv_2[206]) );
  DFFRHQXL conv_2_reg_13__12_ ( .D(n15066), .CK(clk), .RN(rst_n), .Q(
        conv_2[207]) );
  DFFRHQXL conv_2_reg_13__13_ ( .D(n15065), .CK(clk), .RN(rst_n), .Q(
        conv_2[208]) );
  DFFRHQXL conv_2_reg_14__14_ ( .D(n15054), .CK(clk), .RN(rst_n), .Q(
        conv_2[224]) );
  DFFRHQXL conv_2_reg_14__0_ ( .D(n15369), .CK(clk), .RN(rst_n), .Q(
        conv_2[210]) );
  DFFRHQXL conv_2_reg_14__5_ ( .D(n15063), .CK(clk), .RN(rst_n), .Q(
        conv_2[215]) );
  DFFRHQXL conv_2_reg_14__6_ ( .D(n15062), .CK(clk), .RN(rst_n), .Q(
        conv_2[216]) );
  DFFRHQXL conv_2_reg_14__7_ ( .D(n15061), .CK(clk), .RN(rst_n), .Q(
        conv_2[217]) );
  DFFRHQXL conv_2_reg_14__8_ ( .D(n15060), .CK(clk), .RN(rst_n), .Q(
        conv_2[218]) );
  DFFRHQXL conv_2_reg_14__9_ ( .D(n15059), .CK(clk), .RN(rst_n), .Q(
        conv_2[219]) );
  DFFRHQXL conv_2_reg_14__10_ ( .D(n15058), .CK(clk), .RN(rst_n), .Q(
        conv_2[220]) );
  DFFRHQXL conv_2_reg_14__11_ ( .D(n15057), .CK(clk), .RN(rst_n), .Q(
        conv_2[221]) );
  DFFRHQXL conv_2_reg_14__12_ ( .D(n15056), .CK(clk), .RN(rst_n), .Q(
        conv_2[222]) );
  DFFRHQXL conv_2_reg_14__13_ ( .D(n15055), .CK(clk), .RN(rst_n), .Q(
        conv_2[223]) );
  DFFRHQXL conv_2_reg_15__14_ ( .D(n15044), .CK(clk), .RN(rst_n), .Q(
        conv_2[239]) );
  DFFRHQXL conv_2_reg_15__0_ ( .D(n15368), .CK(clk), .RN(rst_n), .Q(
        conv_2[225]) );
  DFFRHQXL conv_2_reg_15__5_ ( .D(n15053), .CK(clk), .RN(rst_n), .Q(
        conv_2[230]) );
  DFFRHQXL conv_2_reg_15__6_ ( .D(n15052), .CK(clk), .RN(rst_n), .Q(
        conv_2[231]) );
  DFFRHQXL conv_2_reg_15__7_ ( .D(n15051), .CK(clk), .RN(rst_n), .Q(
        conv_2[232]) );
  DFFRHQXL conv_2_reg_15__8_ ( .D(n15050), .CK(clk), .RN(rst_n), .Q(
        conv_2[233]) );
  DFFRHQXL conv_2_reg_15__9_ ( .D(n15049), .CK(clk), .RN(rst_n), .Q(
        conv_2[234]) );
  DFFRHQXL conv_2_reg_15__10_ ( .D(n15048), .CK(clk), .RN(rst_n), .Q(
        conv_2[235]) );
  DFFRHQXL conv_2_reg_15__11_ ( .D(n15047), .CK(clk), .RN(rst_n), .Q(
        conv_2[236]) );
  DFFRHQXL conv_2_reg_15__12_ ( .D(n15046), .CK(clk), .RN(rst_n), .Q(
        conv_2[237]) );
  DFFRHQXL conv_2_reg_15__13_ ( .D(n15045), .CK(clk), .RN(rst_n), .Q(
        conv_2[238]) );
  DFFRHQXL conv_2_reg_16__14_ ( .D(n15034), .CK(clk), .RN(rst_n), .Q(
        conv_2[254]) );
  DFFRHQXL conv_2_reg_16__0_ ( .D(n15367), .CK(clk), .RN(rst_n), .Q(
        conv_2[240]) );
  DFFRHQXL conv_2_reg_16__5_ ( .D(n15043), .CK(clk), .RN(rst_n), .Q(
        conv_2[245]) );
  DFFRHQXL conv_2_reg_16__6_ ( .D(n15042), .CK(clk), .RN(rst_n), .Q(
        conv_2[246]) );
  DFFRHQXL conv_2_reg_16__7_ ( .D(n15041), .CK(clk), .RN(rst_n), .Q(
        conv_2[247]) );
  DFFRHQXL conv_2_reg_16__8_ ( .D(n15040), .CK(clk), .RN(rst_n), .Q(
        conv_2[248]) );
  DFFRHQXL conv_2_reg_16__9_ ( .D(n15039), .CK(clk), .RN(rst_n), .Q(
        conv_2[249]) );
  DFFRHQXL conv_2_reg_16__10_ ( .D(n15038), .CK(clk), .RN(rst_n), .Q(
        conv_2[250]) );
  DFFRHQXL conv_2_reg_16__11_ ( .D(n15037), .CK(clk), .RN(rst_n), .Q(
        conv_2[251]) );
  DFFRHQXL conv_2_reg_16__12_ ( .D(n15036), .CK(clk), .RN(rst_n), .Q(
        conv_2[252]) );
  DFFRHQXL conv_2_reg_16__13_ ( .D(n15035), .CK(clk), .RN(rst_n), .Q(
        conv_2[253]) );
  DFFRHQXL conv_2_reg_17__14_ ( .D(n15024), .CK(clk), .RN(rst_n), .Q(
        conv_2[269]) );
  DFFRHQXL conv_2_reg_17__0_ ( .D(n15366), .CK(clk), .RN(rst_n), .Q(
        conv_2[255]) );
  DFFRHQXL conv_2_reg_17__5_ ( .D(n15033), .CK(clk), .RN(rst_n), .Q(
        conv_2[260]) );
  DFFRHQXL conv_2_reg_17__6_ ( .D(n15032), .CK(clk), .RN(rst_n), .Q(
        conv_2[261]) );
  DFFRHQXL conv_2_reg_17__7_ ( .D(n15031), .CK(clk), .RN(rst_n), .Q(
        conv_2[262]) );
  DFFRHQXL conv_2_reg_17__8_ ( .D(n15030), .CK(clk), .RN(rst_n), .Q(
        conv_2[263]) );
  DFFRHQXL conv_2_reg_17__9_ ( .D(n15029), .CK(clk), .RN(rst_n), .Q(
        conv_2[264]) );
  DFFRHQXL conv_2_reg_17__10_ ( .D(n15028), .CK(clk), .RN(rst_n), .Q(
        conv_2[265]) );
  DFFRHQXL conv_2_reg_17__11_ ( .D(n15027), .CK(clk), .RN(rst_n), .Q(
        conv_2[266]) );
  DFFRHQXL conv_2_reg_17__12_ ( .D(n15026), .CK(clk), .RN(rst_n), .Q(
        conv_2[267]) );
  DFFRHQXL conv_2_reg_17__13_ ( .D(n15025), .CK(clk), .RN(rst_n), .Q(
        conv_2[268]) );
  DFFRHQXL conv_2_reg_18__14_ ( .D(n15014), .CK(clk), .RN(rst_n), .Q(
        conv_2[284]) );
  DFFRHQXL conv_2_reg_18__0_ ( .D(n15365), .CK(clk), .RN(rst_n), .Q(
        conv_2[270]) );
  DFFRHQXL conv_2_reg_18__5_ ( .D(n15023), .CK(clk), .RN(rst_n), .Q(
        conv_2[275]) );
  DFFRHQXL conv_2_reg_18__6_ ( .D(n15022), .CK(clk), .RN(rst_n), .Q(
        conv_2[276]) );
  DFFRHQXL conv_2_reg_18__7_ ( .D(n15021), .CK(clk), .RN(rst_n), .Q(
        conv_2[277]) );
  DFFRHQXL conv_2_reg_18__8_ ( .D(n15020), .CK(clk), .RN(rst_n), .Q(
        conv_2[278]) );
  DFFRHQXL conv_2_reg_18__9_ ( .D(n15019), .CK(clk), .RN(rst_n), .Q(
        conv_2[279]) );
  DFFRHQXL conv_2_reg_18__10_ ( .D(n15018), .CK(clk), .RN(rst_n), .Q(
        conv_2[280]) );
  DFFRHQXL conv_2_reg_18__11_ ( .D(n15017), .CK(clk), .RN(rst_n), .Q(
        conv_2[281]) );
  DFFRHQXL conv_2_reg_18__12_ ( .D(n15016), .CK(clk), .RN(rst_n), .Q(
        conv_2[282]) );
  DFFRHQXL conv_2_reg_18__13_ ( .D(n15015), .CK(clk), .RN(rst_n), .Q(
        conv_2[283]) );
  DFFRHQXL conv_2_reg_19__14_ ( .D(n15004), .CK(clk), .RN(rst_n), .Q(
        conv_2[299]) );
  DFFRHQXL conv_2_reg_19__0_ ( .D(n15364), .CK(clk), .RN(rst_n), .Q(
        conv_2[285]) );
  DFFRHQXL conv_2_reg_19__5_ ( .D(n15013), .CK(clk), .RN(rst_n), .Q(
        conv_2[290]) );
  DFFRHQXL conv_2_reg_19__6_ ( .D(n15012), .CK(clk), .RN(rst_n), .Q(
        conv_2[291]) );
  DFFRHQXL conv_2_reg_19__7_ ( .D(n15011), .CK(clk), .RN(rst_n), .Q(
        conv_2[292]) );
  DFFRHQXL conv_2_reg_19__8_ ( .D(n15010), .CK(clk), .RN(rst_n), .Q(
        conv_2[293]) );
  DFFRHQXL conv_2_reg_19__9_ ( .D(n15009), .CK(clk), .RN(rst_n), .Q(
        conv_2[294]) );
  DFFRHQXL conv_2_reg_19__10_ ( .D(n15008), .CK(clk), .RN(rst_n), .Q(
        conv_2[295]) );
  DFFRHQXL conv_2_reg_19__11_ ( .D(n15007), .CK(clk), .RN(rst_n), .Q(
        conv_2[296]) );
  DFFRHQXL conv_2_reg_19__12_ ( .D(n15006), .CK(clk), .RN(rst_n), .Q(
        conv_2[297]) );
  DFFRHQXL conv_2_reg_19__13_ ( .D(n15005), .CK(clk), .RN(rst_n), .Q(
        conv_2[298]) );
  DFFRHQXL conv_2_reg_20__14_ ( .D(n14994), .CK(clk), .RN(rst_n), .Q(
        conv_2[314]) );
  DFFRHQXL conv_2_reg_20__0_ ( .D(n15363), .CK(clk), .RN(rst_n), .Q(
        conv_2[300]) );
  DFFRHQXL conv_2_reg_20__5_ ( .D(n15003), .CK(clk), .RN(rst_n), .Q(
        conv_2[305]) );
  DFFRHQXL conv_2_reg_20__6_ ( .D(n15002), .CK(clk), .RN(rst_n), .Q(
        conv_2[306]) );
  DFFRHQXL conv_2_reg_20__7_ ( .D(n15001), .CK(clk), .RN(rst_n), .Q(
        conv_2[307]) );
  DFFRHQXL conv_2_reg_20__8_ ( .D(n15000), .CK(clk), .RN(rst_n), .Q(
        conv_2[308]) );
  DFFRHQXL conv_2_reg_20__9_ ( .D(n14999), .CK(clk), .RN(rst_n), .Q(
        conv_2[309]) );
  DFFRHQXL conv_2_reg_20__10_ ( .D(n14998), .CK(clk), .RN(rst_n), .Q(
        conv_2[310]) );
  DFFRHQXL conv_2_reg_20__11_ ( .D(n14997), .CK(clk), .RN(rst_n), .Q(
        conv_2[311]) );
  DFFRHQXL conv_2_reg_20__12_ ( .D(n14996), .CK(clk), .RN(rst_n), .Q(
        conv_2[312]) );
  DFFRHQXL conv_2_reg_20__13_ ( .D(n14995), .CK(clk), .RN(rst_n), .Q(
        conv_2[313]) );
  DFFRHQXL conv_2_reg_21__14_ ( .D(n14984), .CK(clk), .RN(rst_n), .Q(
        conv_2[329]) );
  DFFRHQXL conv_2_reg_21__0_ ( .D(n15362), .CK(clk), .RN(rst_n), .Q(
        conv_2[315]) );
  DFFRHQXL conv_2_reg_21__5_ ( .D(n14993), .CK(clk), .RN(rst_n), .Q(
        conv_2[320]) );
  DFFRHQXL conv_2_reg_21__6_ ( .D(n14992), .CK(clk), .RN(rst_n), .Q(
        conv_2[321]) );
  DFFRHQXL conv_2_reg_21__7_ ( .D(n14991), .CK(clk), .RN(rst_n), .Q(
        conv_2[322]) );
  DFFRHQXL conv_2_reg_21__8_ ( .D(n14990), .CK(clk), .RN(rst_n), .Q(
        conv_2[323]) );
  DFFRHQXL conv_2_reg_21__9_ ( .D(n14989), .CK(clk), .RN(rst_n), .Q(
        conv_2[324]) );
  DFFRHQXL conv_2_reg_21__10_ ( .D(n14988), .CK(clk), .RN(rst_n), .Q(
        conv_2[325]) );
  DFFRHQXL conv_2_reg_21__11_ ( .D(n14987), .CK(clk), .RN(rst_n), .Q(
        conv_2[326]) );
  DFFRHQXL conv_2_reg_21__12_ ( .D(n14986), .CK(clk), .RN(rst_n), .Q(
        conv_2[327]) );
  DFFRHQXL conv_2_reg_21__13_ ( .D(n14985), .CK(clk), .RN(rst_n), .Q(
        conv_2[328]) );
  DFFRHQXL conv_2_reg_22__14_ ( .D(n14974), .CK(clk), .RN(rst_n), .Q(
        conv_2[344]) );
  DFFRHQXL conv_2_reg_22__0_ ( .D(n15361), .CK(clk), .RN(rst_n), .Q(
        conv_2[330]) );
  DFFRHQXL conv_2_reg_22__5_ ( .D(n14983), .CK(clk), .RN(rst_n), .Q(
        conv_2[335]) );
  DFFRHQXL conv_2_reg_22__6_ ( .D(n14982), .CK(clk), .RN(rst_n), .Q(
        conv_2[336]) );
  DFFRHQXL conv_2_reg_22__7_ ( .D(n14981), .CK(clk), .RN(rst_n), .Q(
        conv_2[337]) );
  DFFRHQXL conv_2_reg_22__8_ ( .D(n14980), .CK(clk), .RN(rst_n), .Q(
        conv_2[338]) );
  DFFRHQXL conv_2_reg_22__9_ ( .D(n14979), .CK(clk), .RN(rst_n), .Q(
        conv_2[339]) );
  DFFRHQXL conv_2_reg_22__10_ ( .D(n14978), .CK(clk), .RN(rst_n), .Q(
        conv_2[340]) );
  DFFRHQXL conv_2_reg_22__11_ ( .D(n14977), .CK(clk), .RN(rst_n), .Q(
        conv_2[341]) );
  DFFRHQXL conv_2_reg_22__12_ ( .D(n14976), .CK(clk), .RN(rst_n), .Q(
        conv_2[342]) );
  DFFRHQXL conv_2_reg_22__13_ ( .D(n14975), .CK(clk), .RN(rst_n), .Q(
        conv_2[343]) );
  DFFRHQXL conv_2_reg_23__14_ ( .D(n14964), .CK(clk), .RN(rst_n), .Q(
        conv_2[359]) );
  DFFRHQXL conv_2_reg_23__0_ ( .D(n15360), .CK(clk), .RN(rst_n), .Q(
        conv_2[345]) );
  DFFRHQXL conv_2_reg_23__5_ ( .D(n14973), .CK(clk), .RN(rst_n), .Q(
        conv_2[350]) );
  DFFRHQXL conv_2_reg_23__6_ ( .D(n14972), .CK(clk), .RN(rst_n), .Q(
        conv_2[351]) );
  DFFRHQXL conv_2_reg_23__7_ ( .D(n14971), .CK(clk), .RN(rst_n), .Q(
        conv_2[352]) );
  DFFRHQXL conv_2_reg_23__8_ ( .D(n14970), .CK(clk), .RN(rst_n), .Q(
        conv_2[353]) );
  DFFRHQXL conv_2_reg_23__9_ ( .D(n14969), .CK(clk), .RN(rst_n), .Q(
        conv_2[354]) );
  DFFRHQXL conv_2_reg_23__10_ ( .D(n14968), .CK(clk), .RN(rst_n), .Q(
        conv_2[355]) );
  DFFRHQXL conv_2_reg_23__11_ ( .D(n14967), .CK(clk), .RN(rst_n), .Q(
        conv_2[356]) );
  DFFRHQXL conv_2_reg_23__12_ ( .D(n14966), .CK(clk), .RN(rst_n), .Q(
        conv_2[357]) );
  DFFRHQXL conv_2_reg_23__13_ ( .D(n14965), .CK(clk), .RN(rst_n), .Q(
        conv_2[358]) );
  DFFRHQXL conv_2_reg_24__14_ ( .D(n14954), .CK(clk), .RN(rst_n), .Q(
        conv_2[374]) );
  DFFRHQXL conv_2_reg_24__0_ ( .D(n15359), .CK(clk), .RN(rst_n), .Q(
        conv_2[360]) );
  DFFRHQXL conv_2_reg_24__5_ ( .D(n14963), .CK(clk), .RN(rst_n), .Q(
        conv_2[365]) );
  DFFRHQXL conv_2_reg_24__6_ ( .D(n14962), .CK(clk), .RN(rst_n), .Q(
        conv_2[366]) );
  DFFRHQXL conv_2_reg_24__7_ ( .D(n14961), .CK(clk), .RN(rst_n), .Q(
        conv_2[367]) );
  DFFRHQXL conv_2_reg_24__8_ ( .D(n14960), .CK(clk), .RN(rst_n), .Q(
        conv_2[368]) );
  DFFRHQXL conv_2_reg_24__9_ ( .D(n14959), .CK(clk), .RN(rst_n), .Q(
        conv_2[369]) );
  DFFRHQXL conv_2_reg_24__10_ ( .D(n14958), .CK(clk), .RN(rst_n), .Q(
        conv_2[370]) );
  DFFRHQXL conv_2_reg_24__11_ ( .D(n14957), .CK(clk), .RN(rst_n), .Q(
        conv_2[371]) );
  DFFRHQXL conv_2_reg_24__12_ ( .D(n14956), .CK(clk), .RN(rst_n), .Q(
        conv_2[372]) );
  DFFRHQXL conv_2_reg_24__13_ ( .D(n14955), .CK(clk), .RN(rst_n), .Q(
        conv_2[373]) );
  DFFRHQXL conv_2_reg_25__14_ ( .D(n14944), .CK(clk), .RN(rst_n), .Q(
        conv_2[389]) );
  DFFRHQXL conv_2_reg_25__0_ ( .D(n15358), .CK(clk), .RN(rst_n), .Q(
        conv_2[375]) );
  DFFRHQXL conv_2_reg_25__5_ ( .D(n14953), .CK(clk), .RN(rst_n), .Q(
        conv_2[380]) );
  DFFRHQXL conv_2_reg_25__6_ ( .D(n14952), .CK(clk), .RN(rst_n), .Q(
        conv_2[381]) );
  DFFRHQXL conv_2_reg_25__7_ ( .D(n14951), .CK(clk), .RN(rst_n), .Q(
        conv_2[382]) );
  DFFRHQXL conv_2_reg_25__8_ ( .D(n14950), .CK(clk), .RN(rst_n), .Q(
        conv_2[383]) );
  DFFRHQXL conv_2_reg_25__9_ ( .D(n14949), .CK(clk), .RN(rst_n), .Q(
        conv_2[384]) );
  DFFRHQXL conv_2_reg_25__10_ ( .D(n14948), .CK(clk), .RN(rst_n), .Q(
        conv_2[385]) );
  DFFRHQXL conv_2_reg_25__11_ ( .D(n14947), .CK(clk), .RN(rst_n), .Q(
        conv_2[386]) );
  DFFRHQXL conv_2_reg_25__12_ ( .D(n14946), .CK(clk), .RN(rst_n), .Q(
        conv_2[387]) );
  DFFRHQXL conv_2_reg_25__13_ ( .D(n14945), .CK(clk), .RN(rst_n), .Q(
        conv_2[388]) );
  DFFRHQXL conv_2_reg_26__14_ ( .D(n14934), .CK(clk), .RN(rst_n), .Q(
        conv_2[404]) );
  DFFRHQXL conv_2_reg_26__0_ ( .D(n15357), .CK(clk), .RN(rst_n), .Q(
        conv_2[390]) );
  DFFRHQXL conv_2_reg_26__5_ ( .D(n14943), .CK(clk), .RN(rst_n), .Q(
        conv_2[395]) );
  DFFRHQXL conv_2_reg_26__6_ ( .D(n14942), .CK(clk), .RN(rst_n), .Q(
        conv_2[396]) );
  DFFRHQXL conv_2_reg_26__7_ ( .D(n14941), .CK(clk), .RN(rst_n), .Q(
        conv_2[397]) );
  DFFRHQXL conv_2_reg_26__8_ ( .D(n14940), .CK(clk), .RN(rst_n), .Q(
        conv_2[398]) );
  DFFRHQXL conv_2_reg_26__9_ ( .D(n14939), .CK(clk), .RN(rst_n), .Q(
        conv_2[399]) );
  DFFRHQXL conv_2_reg_26__10_ ( .D(n14938), .CK(clk), .RN(rst_n), .Q(
        conv_2[400]) );
  DFFRHQXL conv_2_reg_26__11_ ( .D(n14937), .CK(clk), .RN(rst_n), .Q(
        conv_2[401]) );
  DFFRHQXL conv_2_reg_26__12_ ( .D(n14936), .CK(clk), .RN(rst_n), .Q(
        conv_2[402]) );
  DFFRHQXL conv_2_reg_26__13_ ( .D(n14935), .CK(clk), .RN(rst_n), .Q(
        conv_2[403]) );
  DFFRHQXL conv_2_reg_27__14_ ( .D(n14924), .CK(clk), .RN(rst_n), .Q(
        conv_2[419]) );
  DFFRHQXL conv_2_reg_27__0_ ( .D(n15356), .CK(clk), .RN(rst_n), .Q(
        conv_2[405]) );
  DFFRHQXL conv_2_reg_27__5_ ( .D(n14933), .CK(clk), .RN(rst_n), .Q(
        conv_2[410]) );
  DFFRHQXL conv_2_reg_27__6_ ( .D(n14932), .CK(clk), .RN(rst_n), .Q(
        conv_2[411]) );
  DFFRHQXL conv_2_reg_27__7_ ( .D(n14931), .CK(clk), .RN(rst_n), .Q(
        conv_2[412]) );
  DFFRHQXL conv_2_reg_27__8_ ( .D(n14930), .CK(clk), .RN(rst_n), .Q(
        conv_2[413]) );
  DFFRHQXL conv_2_reg_27__9_ ( .D(n14929), .CK(clk), .RN(rst_n), .Q(
        conv_2[414]) );
  DFFRHQXL conv_2_reg_27__10_ ( .D(n14928), .CK(clk), .RN(rst_n), .Q(
        conv_2[415]) );
  DFFRHQXL conv_2_reg_27__11_ ( .D(n14927), .CK(clk), .RN(rst_n), .Q(
        conv_2[416]) );
  DFFRHQXL conv_2_reg_27__12_ ( .D(n14926), .CK(clk), .RN(rst_n), .Q(
        conv_2[417]) );
  DFFRHQXL conv_2_reg_27__13_ ( .D(n14925), .CK(clk), .RN(rst_n), .Q(
        conv_2[418]) );
  DFFRHQXL conv_2_reg_28__14_ ( .D(n14914), .CK(clk), .RN(rst_n), .Q(
        conv_2[434]) );
  DFFRHQXL conv_2_reg_28__0_ ( .D(n15355), .CK(clk), .RN(rst_n), .Q(
        conv_2[420]) );
  DFFRHQXL conv_2_reg_28__5_ ( .D(n14923), .CK(clk), .RN(rst_n), .Q(
        conv_2[425]) );
  DFFRHQXL conv_2_reg_28__6_ ( .D(n14922), .CK(clk), .RN(rst_n), .Q(
        conv_2[426]) );
  DFFRHQXL conv_2_reg_28__7_ ( .D(n14921), .CK(clk), .RN(rst_n), .Q(
        conv_2[427]) );
  DFFRHQXL conv_2_reg_28__8_ ( .D(n14920), .CK(clk), .RN(rst_n), .Q(
        conv_2[428]) );
  DFFRHQXL conv_2_reg_28__9_ ( .D(n14919), .CK(clk), .RN(rst_n), .Q(
        conv_2[429]) );
  DFFRHQXL conv_2_reg_28__10_ ( .D(n14918), .CK(clk), .RN(rst_n), .Q(
        conv_2[430]) );
  DFFRHQXL conv_2_reg_28__11_ ( .D(n14917), .CK(clk), .RN(rst_n), .Q(
        conv_2[431]) );
  DFFRHQXL conv_2_reg_28__12_ ( .D(n14916), .CK(clk), .RN(rst_n), .Q(
        conv_2[432]) );
  DFFRHQXL conv_2_reg_28__13_ ( .D(n14915), .CK(clk), .RN(rst_n), .Q(
        conv_2[433]) );
  DFFRHQXL conv_2_reg_29__14_ ( .D(n14904), .CK(clk), .RN(rst_n), .Q(
        conv_2[449]) );
  DFFRHQXL conv_2_reg_29__0_ ( .D(n15354), .CK(clk), .RN(rst_n), .Q(
        conv_2[435]) );
  DFFRHQXL conv_2_reg_29__5_ ( .D(n14913), .CK(clk), .RN(rst_n), .Q(
        conv_2[440]) );
  DFFRHQXL conv_2_reg_29__6_ ( .D(n14912), .CK(clk), .RN(rst_n), .Q(
        conv_2[441]) );
  DFFRHQXL conv_2_reg_29__7_ ( .D(n14911), .CK(clk), .RN(rst_n), .Q(
        conv_2[442]) );
  DFFRHQXL conv_2_reg_29__8_ ( .D(n14910), .CK(clk), .RN(rst_n), .Q(
        conv_2[443]) );
  DFFRHQXL conv_2_reg_29__9_ ( .D(n14909), .CK(clk), .RN(rst_n), .Q(
        conv_2[444]) );
  DFFRHQXL conv_2_reg_29__10_ ( .D(n14908), .CK(clk), .RN(rst_n), .Q(
        conv_2[445]) );
  DFFRHQXL conv_2_reg_29__11_ ( .D(n14907), .CK(clk), .RN(rst_n), .Q(
        conv_2[446]) );
  DFFRHQXL conv_2_reg_29__12_ ( .D(n14906), .CK(clk), .RN(rst_n), .Q(
        conv_2[447]) );
  DFFRHQXL conv_2_reg_29__13_ ( .D(n14905), .CK(clk), .RN(rst_n), .Q(
        conv_2[448]) );
  DFFRHQXL conv_2_reg_30__14_ ( .D(n14894), .CK(clk), .RN(rst_n), .Q(
        conv_2[464]) );
  DFFRHQXL conv_2_reg_30__0_ ( .D(n15353), .CK(clk), .RN(rst_n), .Q(
        conv_2[450]) );
  DFFRHQXL conv_2_reg_30__5_ ( .D(n14903), .CK(clk), .RN(rst_n), .Q(
        conv_2[455]) );
  DFFRHQXL conv_2_reg_30__6_ ( .D(n14902), .CK(clk), .RN(rst_n), .Q(
        conv_2[456]) );
  DFFRHQXL conv_2_reg_30__7_ ( .D(n14901), .CK(clk), .RN(rst_n), .Q(
        conv_2[457]) );
  DFFRHQXL conv_2_reg_30__8_ ( .D(n14900), .CK(clk), .RN(rst_n), .Q(
        conv_2[458]) );
  DFFRHQXL conv_2_reg_30__9_ ( .D(n14899), .CK(clk), .RN(rst_n), .Q(
        conv_2[459]) );
  DFFRHQXL conv_2_reg_30__10_ ( .D(n14898), .CK(clk), .RN(rst_n), .Q(
        conv_2[460]) );
  DFFRHQXL conv_2_reg_30__11_ ( .D(n14897), .CK(clk), .RN(rst_n), .Q(
        conv_2[461]) );
  DFFRHQXL conv_2_reg_30__12_ ( .D(n14896), .CK(clk), .RN(rst_n), .Q(
        conv_2[462]) );
  DFFRHQXL conv_2_reg_30__13_ ( .D(n14895), .CK(clk), .RN(rst_n), .Q(
        conv_2[463]) );
  DFFRHQXL conv_2_reg_31__14_ ( .D(n14884), .CK(clk), .RN(rst_n), .Q(
        conv_2[479]) );
  DFFRHQXL conv_2_reg_31__0_ ( .D(n15352), .CK(clk), .RN(rst_n), .Q(
        conv_2[465]) );
  DFFRHQXL conv_2_reg_31__5_ ( .D(n14893), .CK(clk), .RN(rst_n), .Q(
        conv_2[470]) );
  DFFRHQXL conv_2_reg_31__6_ ( .D(n14892), .CK(clk), .RN(rst_n), .Q(
        conv_2[471]) );
  DFFRHQXL conv_2_reg_31__7_ ( .D(n14891), .CK(clk), .RN(rst_n), .Q(
        conv_2[472]) );
  DFFRHQXL conv_2_reg_31__8_ ( .D(n14890), .CK(clk), .RN(rst_n), .Q(
        conv_2[473]) );
  DFFRHQXL conv_2_reg_31__9_ ( .D(n14889), .CK(clk), .RN(rst_n), .Q(
        conv_2[474]) );
  DFFRHQXL conv_2_reg_31__10_ ( .D(n14888), .CK(clk), .RN(rst_n), .Q(
        conv_2[475]) );
  DFFRHQXL conv_2_reg_31__11_ ( .D(n14887), .CK(clk), .RN(rst_n), .Q(
        conv_2[476]) );
  DFFRHQXL conv_2_reg_31__12_ ( .D(n14886), .CK(clk), .RN(rst_n), .Q(
        conv_2[477]) );
  DFFRHQXL conv_2_reg_31__13_ ( .D(n14885), .CK(clk), .RN(rst_n), .Q(
        conv_2[478]) );
  DFFRHQXL conv_2_reg_32__14_ ( .D(n14874), .CK(clk), .RN(rst_n), .Q(
        conv_2[494]) );
  DFFRHQXL conv_2_reg_32__0_ ( .D(n15351), .CK(clk), .RN(rst_n), .Q(
        conv_2[480]) );
  DFFRHQXL conv_2_reg_32__5_ ( .D(n14883), .CK(clk), .RN(rst_n), .Q(
        conv_2[485]) );
  DFFRHQXL conv_2_reg_32__6_ ( .D(n14882), .CK(clk), .RN(rst_n), .Q(
        conv_2[486]) );
  DFFRHQXL conv_2_reg_32__7_ ( .D(n14881), .CK(clk), .RN(rst_n), .Q(
        conv_2[487]) );
  DFFRHQXL conv_2_reg_32__8_ ( .D(n14880), .CK(clk), .RN(rst_n), .Q(
        conv_2[488]) );
  DFFRHQXL conv_2_reg_32__9_ ( .D(n14879), .CK(clk), .RN(rst_n), .Q(
        conv_2[489]) );
  DFFRHQXL conv_2_reg_32__10_ ( .D(n14878), .CK(clk), .RN(rst_n), .Q(
        conv_2[490]) );
  DFFRHQXL conv_2_reg_32__11_ ( .D(n14877), .CK(clk), .RN(rst_n), .Q(
        conv_2[491]) );
  DFFRHQXL conv_2_reg_32__12_ ( .D(n14876), .CK(clk), .RN(rst_n), .Q(
        conv_2[492]) );
  DFFRHQXL conv_2_reg_32__13_ ( .D(n14875), .CK(clk), .RN(rst_n), .Q(
        conv_2[493]) );
  DFFRHQXL conv_2_reg_33__14_ ( .D(n14864), .CK(clk), .RN(rst_n), .Q(
        conv_2[509]) );
  DFFRHQXL conv_2_reg_33__0_ ( .D(n15350), .CK(clk), .RN(rst_n), .Q(
        conv_2[495]) );
  DFFRHQXL conv_2_reg_33__5_ ( .D(n14873), .CK(clk), .RN(rst_n), .Q(
        conv_2[500]) );
  DFFRHQXL conv_2_reg_33__6_ ( .D(n14872), .CK(clk), .RN(rst_n), .Q(
        conv_2[501]) );
  DFFRHQXL conv_2_reg_33__7_ ( .D(n14871), .CK(clk), .RN(rst_n), .Q(
        conv_2[502]) );
  DFFRHQXL conv_2_reg_33__8_ ( .D(n14870), .CK(clk), .RN(rst_n), .Q(
        conv_2[503]) );
  DFFRHQXL conv_2_reg_33__9_ ( .D(n14869), .CK(clk), .RN(rst_n), .Q(
        conv_2[504]) );
  DFFRHQXL conv_2_reg_33__10_ ( .D(n14868), .CK(clk), .RN(rst_n), .Q(
        conv_2[505]) );
  DFFRHQXL conv_2_reg_33__11_ ( .D(n14867), .CK(clk), .RN(rst_n), .Q(
        conv_2[506]) );
  DFFRHQXL conv_2_reg_33__12_ ( .D(n14866), .CK(clk), .RN(rst_n), .Q(
        conv_2[507]) );
  DFFRHQXL conv_2_reg_33__13_ ( .D(n14865), .CK(clk), .RN(rst_n), .Q(
        conv_2[508]) );
  DFFRHQXL conv_2_reg_34__14_ ( .D(n14854), .CK(clk), .RN(rst_n), .Q(
        conv_2[524]) );
  DFFRHQXL conv_2_reg_34__0_ ( .D(n15349), .CK(clk), .RN(rst_n), .Q(
        conv_2[510]) );
  DFFRHQXL conv_2_reg_34__5_ ( .D(n14863), .CK(clk), .RN(rst_n), .Q(
        conv_2[515]) );
  DFFRHQXL conv_2_reg_34__6_ ( .D(n14862), .CK(clk), .RN(rst_n), .Q(
        conv_2[516]) );
  DFFRHQXL conv_2_reg_34__7_ ( .D(n14861), .CK(clk), .RN(rst_n), .Q(
        conv_2[517]) );
  DFFRHQXL conv_2_reg_34__8_ ( .D(n14860), .CK(clk), .RN(rst_n), .Q(
        conv_2[518]) );
  DFFRHQXL conv_2_reg_34__9_ ( .D(n14859), .CK(clk), .RN(rst_n), .Q(
        conv_2[519]) );
  DFFRHQXL conv_2_reg_34__10_ ( .D(n14858), .CK(clk), .RN(rst_n), .Q(
        conv_2[520]) );
  DFFRHQXL conv_2_reg_34__11_ ( .D(n14857), .CK(clk), .RN(rst_n), .Q(
        conv_2[521]) );
  DFFRHQXL conv_2_reg_34__12_ ( .D(n14856), .CK(clk), .RN(rst_n), .Q(
        conv_2[522]) );
  DFFRHQXL conv_2_reg_34__13_ ( .D(n14855), .CK(clk), .RN(rst_n), .Q(
        conv_2[523]) );
  DFFRHQXL conv_2_reg_35__14_ ( .D(n14844), .CK(clk), .RN(rst_n), .Q(
        conv_2[539]) );
  DFFRHQXL conv_2_reg_35__0_ ( .D(n15348), .CK(clk), .RN(rst_n), .Q(
        conv_2[525]) );
  DFFRHQXL pool_reg_15__0_ ( .D(N29291), .CK(clk), .RN(rst_n), .Q(pool[75]) );
  DFFRHQXL pool_reg_17__0_ ( .D(N29301), .CK(clk), .RN(rst_n), .Q(pool[85]) );
  DFFRHQXL pool_reg_12__0_ ( .D(N29276), .CK(clk), .RN(rst_n), .Q(pool[60]) );
  DFFRHQXL pool_reg_11__0_ ( .D(N29271), .CK(clk), .RN(rst_n), .Q(pool[55]) );
  DFFRHQXL pool_reg_14__0_ ( .D(N29286), .CK(clk), .RN(rst_n), .Q(pool[70]) );
  DFFRHQXL pool_reg_9__0_ ( .D(N29261), .CK(clk), .RN(rst_n), .Q(pool[45]) );
  DFFRHQXL pool_reg_10__0_ ( .D(N29266), .CK(clk), .RN(rst_n), .Q(pool[50]) );
  DFFRHQXL pool_reg_16__0_ ( .D(N29296), .CK(clk), .RN(rst_n), .Q(pool[80]) );
  DFFRHQXL pool_reg_13__0_ ( .D(N29281), .CK(clk), .RN(rst_n), .Q(pool[65]) );
  DFFRHQXL conv_2_reg_35__5_ ( .D(n14853), .CK(clk), .RN(rst_n), .Q(
        conv_2[530]) );
  DFFRHQXL conv_2_reg_35__6_ ( .D(n14852), .CK(clk), .RN(rst_n), .Q(
        conv_2[531]) );
  DFFRHQXL conv_2_reg_35__7_ ( .D(n14851), .CK(clk), .RN(rst_n), .Q(
        conv_2[532]) );
  DFFRHQXL conv_2_reg_35__8_ ( .D(n14850), .CK(clk), .RN(rst_n), .Q(
        conv_2[533]) );
  DFFRHQXL conv_2_reg_35__9_ ( .D(n14849), .CK(clk), .RN(rst_n), .Q(
        conv_2[534]) );
  DFFRHQXL conv_2_reg_35__10_ ( .D(n14848), .CK(clk), .RN(rst_n), .Q(
        conv_2[535]) );
  DFFRHQXL conv_2_reg_35__11_ ( .D(n14847), .CK(clk), .RN(rst_n), .Q(
        conv_2[536]) );
  DFFRHQXL conv_2_reg_35__12_ ( .D(n14846), .CK(clk), .RN(rst_n), .Q(
        conv_2[537]) );
  DFFRHQXL conv_2_reg_35__13_ ( .D(n14845), .CK(clk), .RN(rst_n), .Q(
        conv_2[538]) );
  DFFRHQXL filter_1_bias_reg_5_ ( .D(n14730), .CK(clk), .RN(rst_n), .Q(
        filter_1_bias[5]) );
  DFFRHQXL conv_1_reg_0__14_ ( .D(n16449), .CK(clk), .RN(rst_n), .Q(conv_1[14]) );
  DFFRHQXL conv_1_reg_0__0_ ( .D(n16463), .CK(clk), .RN(rst_n), .Q(conv_1[0])
         );
  DFFRHQXL conv_1_reg_0__5_ ( .D(n16458), .CK(clk), .RN(rst_n), .Q(conv_1[5])
         );
  DFFRHQXL conv_1_reg_0__6_ ( .D(n16457), .CK(clk), .RN(rst_n), .Q(conv_1[6])
         );
  DFFRHQXL conv_1_reg_0__7_ ( .D(n16456), .CK(clk), .RN(rst_n), .Q(conv_1[7])
         );
  DFFRHQXL conv_1_reg_0__8_ ( .D(n16455), .CK(clk), .RN(rst_n), .Q(conv_1[8])
         );
  DFFRHQXL conv_1_reg_0__9_ ( .D(n16454), .CK(clk), .RN(rst_n), .Q(conv_1[9])
         );
  DFFRHQXL conv_1_reg_0__10_ ( .D(n16453), .CK(clk), .RN(rst_n), .Q(conv_1[10]) );
  DFFRHQXL conv_1_reg_0__11_ ( .D(n16452), .CK(clk), .RN(rst_n), .Q(conv_1[11]) );
  DFFRHQXL conv_1_reg_0__12_ ( .D(n16451), .CK(clk), .RN(rst_n), .Q(conv_1[12]) );
  DFFRHQXL conv_1_reg_0__13_ ( .D(n16450), .CK(clk), .RN(rst_n), .Q(conv_1[13]) );
  DFFRHQXL conv_1_reg_1__14_ ( .D(n16434), .CK(clk), .RN(rst_n), .Q(conv_1[29]) );
  DFFRHQXL conv_1_reg_1__0_ ( .D(n16448), .CK(clk), .RN(rst_n), .Q(conv_1[15])
         );
  DFFRHQXL conv_1_reg_1__5_ ( .D(n16443), .CK(clk), .RN(rst_n), .Q(conv_1[20])
         );
  DFFRHQXL conv_1_reg_1__6_ ( .D(n16442), .CK(clk), .RN(rst_n), .Q(conv_1[21])
         );
  DFFRHQXL conv_1_reg_1__7_ ( .D(n16441), .CK(clk), .RN(rst_n), .Q(conv_1[22])
         );
  DFFRHQXL conv_1_reg_1__8_ ( .D(n16440), .CK(clk), .RN(rst_n), .Q(conv_1[23])
         );
  DFFRHQXL conv_1_reg_1__9_ ( .D(n16439), .CK(clk), .RN(rst_n), .Q(conv_1[24])
         );
  DFFRHQXL conv_1_reg_1__10_ ( .D(n16438), .CK(clk), .RN(rst_n), .Q(conv_1[25]) );
  DFFRHQXL conv_1_reg_1__11_ ( .D(n16437), .CK(clk), .RN(rst_n), .Q(conv_1[26]) );
  DFFRHQXL conv_1_reg_1__12_ ( .D(n16436), .CK(clk), .RN(rst_n), .Q(conv_1[27]) );
  DFFRHQXL conv_1_reg_1__13_ ( .D(n16435), .CK(clk), .RN(rst_n), .Q(conv_1[28]) );
  DFFRHQXL conv_1_reg_2__14_ ( .D(n16419), .CK(clk), .RN(rst_n), .Q(conv_1[44]) );
  DFFRHQXL conv_1_reg_2__0_ ( .D(n16433), .CK(clk), .RN(rst_n), .Q(conv_1[30])
         );
  DFFRHQXL conv_1_reg_2__5_ ( .D(n16428), .CK(clk), .RN(rst_n), .Q(conv_1[35])
         );
  DFFRHQXL conv_1_reg_2__6_ ( .D(n16427), .CK(clk), .RN(rst_n), .Q(conv_1[36])
         );
  DFFRHQXL conv_1_reg_2__7_ ( .D(n16426), .CK(clk), .RN(rst_n), .Q(conv_1[37])
         );
  DFFRHQXL conv_1_reg_2__8_ ( .D(n16425), .CK(clk), .RN(rst_n), .Q(conv_1[38])
         );
  DFFRHQXL conv_1_reg_2__9_ ( .D(n16424), .CK(clk), .RN(rst_n), .Q(conv_1[39])
         );
  DFFRHQXL conv_1_reg_2__10_ ( .D(n16423), .CK(clk), .RN(rst_n), .Q(conv_1[40]) );
  DFFRHQXL conv_1_reg_2__11_ ( .D(n16422), .CK(clk), .RN(rst_n), .Q(conv_1[41]) );
  DFFRHQXL conv_1_reg_2__12_ ( .D(n16421), .CK(clk), .RN(rst_n), .Q(conv_1[42]) );
  DFFRHQXL conv_1_reg_2__13_ ( .D(n16420), .CK(clk), .RN(rst_n), .Q(conv_1[43]) );
  DFFRHQXL conv_1_reg_3__14_ ( .D(n16404), .CK(clk), .RN(rst_n), .Q(conv_1[59]) );
  DFFRHQXL conv_1_reg_3__0_ ( .D(n16418), .CK(clk), .RN(rst_n), .Q(conv_1[45])
         );
  DFFRHQXL conv_1_reg_3__5_ ( .D(n16413), .CK(clk), .RN(rst_n), .Q(conv_1[50])
         );
  DFFRHQXL conv_1_reg_3__6_ ( .D(n16412), .CK(clk), .RN(rst_n), .Q(conv_1[51])
         );
  DFFRHQXL conv_1_reg_3__7_ ( .D(n16411), .CK(clk), .RN(rst_n), .Q(conv_1[52])
         );
  DFFRHQXL conv_1_reg_3__8_ ( .D(n16410), .CK(clk), .RN(rst_n), .Q(conv_1[53])
         );
  DFFRHQXL conv_1_reg_3__9_ ( .D(n16409), .CK(clk), .RN(rst_n), .Q(conv_1[54])
         );
  DFFRHQXL conv_1_reg_3__10_ ( .D(n16408), .CK(clk), .RN(rst_n), .Q(conv_1[55]) );
  DFFRHQXL conv_1_reg_3__11_ ( .D(n16407), .CK(clk), .RN(rst_n), .Q(conv_1[56]) );
  DFFRHQXL conv_1_reg_3__12_ ( .D(n16406), .CK(clk), .RN(rst_n), .Q(conv_1[57]) );
  DFFRHQXL conv_1_reg_3__13_ ( .D(n16405), .CK(clk), .RN(rst_n), .Q(conv_1[58]) );
  DFFRHQXL conv_1_reg_4__14_ ( .D(n16389), .CK(clk), .RN(rst_n), .Q(conv_1[74]) );
  DFFRHQXL conv_1_reg_4__0_ ( .D(n16403), .CK(clk), .RN(rst_n), .Q(conv_1[60])
         );
  DFFRHQXL conv_1_reg_4__5_ ( .D(n16398), .CK(clk), .RN(rst_n), .Q(conv_1[65])
         );
  DFFRHQXL conv_1_reg_4__6_ ( .D(n16397), .CK(clk), .RN(rst_n), .Q(conv_1[66])
         );
  DFFRHQXL conv_1_reg_4__7_ ( .D(n16396), .CK(clk), .RN(rst_n), .Q(conv_1[67])
         );
  DFFRHQXL conv_1_reg_4__8_ ( .D(n16395), .CK(clk), .RN(rst_n), .Q(conv_1[68])
         );
  DFFRHQXL conv_1_reg_4__9_ ( .D(n16394), .CK(clk), .RN(rst_n), .Q(conv_1[69])
         );
  DFFRHQXL conv_1_reg_4__10_ ( .D(n16393), .CK(clk), .RN(rst_n), .Q(conv_1[70]) );
  DFFRHQXL conv_1_reg_4__11_ ( .D(n16392), .CK(clk), .RN(rst_n), .Q(conv_1[71]) );
  DFFRHQXL conv_1_reg_4__12_ ( .D(n16391), .CK(clk), .RN(rst_n), .Q(conv_1[72]) );
  DFFRHQXL conv_1_reg_4__13_ ( .D(n16390), .CK(clk), .RN(rst_n), .Q(conv_1[73]) );
  DFFRHQXL conv_1_reg_5__14_ ( .D(n16374), .CK(clk), .RN(rst_n), .Q(conv_1[89]) );
  DFFRHQXL conv_1_reg_5__0_ ( .D(n16388), .CK(clk), .RN(rst_n), .Q(conv_1[75])
         );
  DFFRHQXL conv_1_reg_5__5_ ( .D(n16383), .CK(clk), .RN(rst_n), .Q(conv_1[80])
         );
  DFFRHQXL conv_1_reg_5__6_ ( .D(n16382), .CK(clk), .RN(rst_n), .Q(conv_1[81])
         );
  DFFRHQXL conv_1_reg_5__7_ ( .D(n16381), .CK(clk), .RN(rst_n), .Q(conv_1[82])
         );
  DFFRHQXL conv_1_reg_5__8_ ( .D(n16380), .CK(clk), .RN(rst_n), .Q(conv_1[83])
         );
  DFFRHQXL conv_1_reg_5__9_ ( .D(n16379), .CK(clk), .RN(rst_n), .Q(conv_1[84])
         );
  DFFRHQXL conv_1_reg_5__10_ ( .D(n16378), .CK(clk), .RN(rst_n), .Q(conv_1[85]) );
  DFFRHQXL conv_1_reg_5__11_ ( .D(n16377), .CK(clk), .RN(rst_n), .Q(conv_1[86]) );
  DFFRHQXL conv_1_reg_5__12_ ( .D(n16376), .CK(clk), .RN(rst_n), .Q(conv_1[87]) );
  DFFRHQXL conv_1_reg_5__13_ ( .D(n16375), .CK(clk), .RN(rst_n), .Q(conv_1[88]) );
  DFFRHQXL conv_1_reg_6__14_ ( .D(n16359), .CK(clk), .RN(rst_n), .Q(
        conv_1[104]) );
  DFFRHQXL conv_1_reg_6__0_ ( .D(n16373), .CK(clk), .RN(rst_n), .Q(conv_1[90])
         );
  DFFRHQXL conv_1_reg_6__5_ ( .D(n16368), .CK(clk), .RN(rst_n), .Q(conv_1[95])
         );
  DFFRHQXL conv_1_reg_6__6_ ( .D(n16367), .CK(clk), .RN(rst_n), .Q(conv_1[96])
         );
  DFFRHQXL conv_1_reg_6__7_ ( .D(n16366), .CK(clk), .RN(rst_n), .Q(conv_1[97])
         );
  DFFRHQXL conv_1_reg_6__8_ ( .D(n16365), .CK(clk), .RN(rst_n), .Q(conv_1[98])
         );
  DFFRHQXL conv_1_reg_6__9_ ( .D(n16364), .CK(clk), .RN(rst_n), .Q(conv_1[99])
         );
  DFFRHQXL conv_1_reg_6__10_ ( .D(n16363), .CK(clk), .RN(rst_n), .Q(
        conv_1[100]) );
  DFFRHQXL conv_1_reg_6__11_ ( .D(n16362), .CK(clk), .RN(rst_n), .Q(
        conv_1[101]) );
  DFFRHQXL conv_1_reg_6__12_ ( .D(n16361), .CK(clk), .RN(rst_n), .Q(
        conv_1[102]) );
  DFFRHQXL conv_1_reg_6__13_ ( .D(n16360), .CK(clk), .RN(rst_n), .Q(
        conv_1[103]) );
  DFFRHQXL conv_1_reg_7__14_ ( .D(n16344), .CK(clk), .RN(rst_n), .Q(
        conv_1[119]) );
  DFFRHQXL conv_1_reg_7__0_ ( .D(n16358), .CK(clk), .RN(rst_n), .Q(conv_1[105]) );
  DFFRHQXL conv_1_reg_7__5_ ( .D(n16353), .CK(clk), .RN(rst_n), .Q(conv_1[110]) );
  DFFRHQXL conv_1_reg_7__6_ ( .D(n16352), .CK(clk), .RN(rst_n), .Q(conv_1[111]) );
  DFFRHQXL conv_1_reg_7__7_ ( .D(n16351), .CK(clk), .RN(rst_n), .Q(conv_1[112]) );
  DFFRHQXL conv_1_reg_7__8_ ( .D(n16350), .CK(clk), .RN(rst_n), .Q(conv_1[113]) );
  DFFRHQXL conv_1_reg_7__9_ ( .D(n16349), .CK(clk), .RN(rst_n), .Q(conv_1[114]) );
  DFFRHQXL conv_1_reg_7__10_ ( .D(n16348), .CK(clk), .RN(rst_n), .Q(
        conv_1[115]) );
  DFFRHQXL conv_1_reg_7__11_ ( .D(n16347), .CK(clk), .RN(rst_n), .Q(
        conv_1[116]) );
  DFFRHQXL conv_1_reg_7__12_ ( .D(n16346), .CK(clk), .RN(rst_n), .Q(
        conv_1[117]) );
  DFFRHQXL conv_1_reg_7__13_ ( .D(n16345), .CK(clk), .RN(rst_n), .Q(
        conv_1[118]) );
  DFFRHQXL conv_1_reg_8__14_ ( .D(n16329), .CK(clk), .RN(rst_n), .Q(
        conv_1[134]) );
  DFFRHQXL conv_1_reg_8__0_ ( .D(n16343), .CK(clk), .RN(rst_n), .Q(conv_1[120]) );
  DFFRHQXL conv_1_reg_8__5_ ( .D(n16338), .CK(clk), .RN(rst_n), .Q(conv_1[125]) );
  DFFRHQXL conv_1_reg_8__6_ ( .D(n16337), .CK(clk), .RN(rst_n), .Q(conv_1[126]) );
  DFFRHQXL conv_1_reg_8__7_ ( .D(n16336), .CK(clk), .RN(rst_n), .Q(conv_1[127]) );
  DFFRHQXL conv_1_reg_8__8_ ( .D(n16335), .CK(clk), .RN(rst_n), .Q(conv_1[128]) );
  DFFRHQXL conv_1_reg_8__9_ ( .D(n16334), .CK(clk), .RN(rst_n), .Q(conv_1[129]) );
  DFFRHQXL conv_1_reg_8__10_ ( .D(n16333), .CK(clk), .RN(rst_n), .Q(
        conv_1[130]) );
  DFFRHQXL conv_1_reg_8__11_ ( .D(n16332), .CK(clk), .RN(rst_n), .Q(
        conv_1[131]) );
  DFFRHQXL conv_1_reg_8__12_ ( .D(n16331), .CK(clk), .RN(rst_n), .Q(
        conv_1[132]) );
  DFFRHQXL conv_1_reg_8__13_ ( .D(n16330), .CK(clk), .RN(rst_n), .Q(
        conv_1[133]) );
  DFFRHQXL conv_1_reg_9__14_ ( .D(n16314), .CK(clk), .RN(rst_n), .Q(
        conv_1[149]) );
  DFFRHQXL conv_1_reg_9__0_ ( .D(n16328), .CK(clk), .RN(rst_n), .Q(conv_1[135]) );
  DFFRHQXL conv_1_reg_9__5_ ( .D(n16323), .CK(clk), .RN(rst_n), .Q(conv_1[140]) );
  DFFRHQXL conv_1_reg_9__6_ ( .D(n16322), .CK(clk), .RN(rst_n), .Q(conv_1[141]) );
  DFFRHQXL conv_1_reg_9__7_ ( .D(n16321), .CK(clk), .RN(rst_n), .Q(conv_1[142]) );
  DFFRHQXL conv_1_reg_9__8_ ( .D(n16320), .CK(clk), .RN(rst_n), .Q(conv_1[143]) );
  DFFRHQXL conv_1_reg_9__9_ ( .D(n16319), .CK(clk), .RN(rst_n), .Q(conv_1[144]) );
  DFFRHQXL conv_1_reg_9__10_ ( .D(n16318), .CK(clk), .RN(rst_n), .Q(
        conv_1[145]) );
  DFFRHQXL conv_1_reg_9__11_ ( .D(n16317), .CK(clk), .RN(rst_n), .Q(
        conv_1[146]) );
  DFFRHQXL conv_1_reg_9__12_ ( .D(n16316), .CK(clk), .RN(rst_n), .Q(
        conv_1[147]) );
  DFFRHQXL conv_1_reg_9__13_ ( .D(n16315), .CK(clk), .RN(rst_n), .Q(
        conv_1[148]) );
  DFFRHQXL conv_1_reg_10__14_ ( .D(n16299), .CK(clk), .RN(rst_n), .Q(
        conv_1[164]) );
  DFFRHQXL conv_1_reg_10__0_ ( .D(n16313), .CK(clk), .RN(rst_n), .Q(
        conv_1[150]) );
  DFFRHQXL conv_1_reg_10__5_ ( .D(n16308), .CK(clk), .RN(rst_n), .Q(
        conv_1[155]) );
  DFFRHQXL conv_1_reg_10__6_ ( .D(n16307), .CK(clk), .RN(rst_n), .Q(
        conv_1[156]) );
  DFFRHQXL conv_1_reg_10__7_ ( .D(n16306), .CK(clk), .RN(rst_n), .Q(
        conv_1[157]) );
  DFFRHQXL conv_1_reg_10__8_ ( .D(n16305), .CK(clk), .RN(rst_n), .Q(
        conv_1[158]) );
  DFFRHQXL conv_1_reg_10__9_ ( .D(n16304), .CK(clk), .RN(rst_n), .Q(
        conv_1[159]) );
  DFFRHQXL conv_1_reg_10__10_ ( .D(n16303), .CK(clk), .RN(rst_n), .Q(
        conv_1[160]) );
  DFFRHQXL conv_1_reg_10__11_ ( .D(n16302), .CK(clk), .RN(rst_n), .Q(
        conv_1[161]) );
  DFFRHQXL conv_1_reg_10__12_ ( .D(n16301), .CK(clk), .RN(rst_n), .Q(
        conv_1[162]) );
  DFFRHQXL conv_1_reg_10__13_ ( .D(n16300), .CK(clk), .RN(rst_n), .Q(
        conv_1[163]) );
  DFFRHQXL conv_1_reg_11__14_ ( .D(n16284), .CK(clk), .RN(rst_n), .Q(
        conv_1[179]) );
  DFFRHQXL conv_1_reg_11__0_ ( .D(n16298), .CK(clk), .RN(rst_n), .Q(
        conv_1[165]) );
  DFFRHQXL conv_1_reg_11__5_ ( .D(n16293), .CK(clk), .RN(rst_n), .Q(
        conv_1[170]) );
  DFFRHQXL conv_1_reg_11__6_ ( .D(n16292), .CK(clk), .RN(rst_n), .Q(
        conv_1[171]) );
  DFFRHQXL conv_1_reg_11__7_ ( .D(n16291), .CK(clk), .RN(rst_n), .Q(
        conv_1[172]) );
  DFFRHQXL conv_1_reg_11__8_ ( .D(n16290), .CK(clk), .RN(rst_n), .Q(
        conv_1[173]) );
  DFFRHQXL conv_1_reg_11__9_ ( .D(n16289), .CK(clk), .RN(rst_n), .Q(
        conv_1[174]) );
  DFFRHQXL conv_1_reg_11__10_ ( .D(n16288), .CK(clk), .RN(rst_n), .Q(
        conv_1[175]) );
  DFFRHQXL conv_1_reg_11__11_ ( .D(n16287), .CK(clk), .RN(rst_n), .Q(
        conv_1[176]) );
  DFFRHQXL conv_1_reg_11__12_ ( .D(n16286), .CK(clk), .RN(rst_n), .Q(
        conv_1[177]) );
  DFFRHQXL conv_1_reg_11__13_ ( .D(n16285), .CK(clk), .RN(rst_n), .Q(
        conv_1[178]) );
  DFFRHQXL conv_1_reg_12__14_ ( .D(n16269), .CK(clk), .RN(rst_n), .Q(
        conv_1[194]) );
  DFFRHQXL conv_1_reg_12__0_ ( .D(n16283), .CK(clk), .RN(rst_n), .Q(
        conv_1[180]) );
  DFFRHQXL conv_1_reg_12__5_ ( .D(n16278), .CK(clk), .RN(rst_n), .Q(
        conv_1[185]) );
  DFFRHQXL conv_1_reg_12__6_ ( .D(n16277), .CK(clk), .RN(rst_n), .Q(
        conv_1[186]) );
  DFFRHQXL conv_1_reg_12__7_ ( .D(n16276), .CK(clk), .RN(rst_n), .Q(
        conv_1[187]) );
  DFFRHQXL conv_1_reg_12__8_ ( .D(n16275), .CK(clk), .RN(rst_n), .Q(
        conv_1[188]) );
  DFFRHQXL conv_1_reg_12__9_ ( .D(n16274), .CK(clk), .RN(rst_n), .Q(
        conv_1[189]) );
  DFFRHQXL conv_1_reg_12__10_ ( .D(n16273), .CK(clk), .RN(rst_n), .Q(
        conv_1[190]) );
  DFFRHQXL conv_1_reg_12__11_ ( .D(n16272), .CK(clk), .RN(rst_n), .Q(
        conv_1[191]) );
  DFFRHQXL conv_1_reg_12__12_ ( .D(n16271), .CK(clk), .RN(rst_n), .Q(
        conv_1[192]) );
  DFFRHQXL conv_1_reg_12__13_ ( .D(n16270), .CK(clk), .RN(rst_n), .Q(
        conv_1[193]) );
  DFFRHQXL conv_1_reg_13__14_ ( .D(n16254), .CK(clk), .RN(rst_n), .Q(
        conv_1[209]) );
  DFFRHQXL conv_1_reg_13__0_ ( .D(n16268), .CK(clk), .RN(rst_n), .Q(
        conv_1[195]) );
  DFFRHQXL conv_1_reg_13__5_ ( .D(n16263), .CK(clk), .RN(rst_n), .Q(
        conv_1[200]) );
  DFFRHQXL conv_1_reg_13__6_ ( .D(n16262), .CK(clk), .RN(rst_n), .Q(
        conv_1[201]) );
  DFFRHQXL conv_1_reg_13__7_ ( .D(n16261), .CK(clk), .RN(rst_n), .Q(
        conv_1[202]) );
  DFFRHQXL conv_1_reg_13__8_ ( .D(n16260), .CK(clk), .RN(rst_n), .Q(
        conv_1[203]) );
  DFFRHQXL conv_1_reg_13__9_ ( .D(n16259), .CK(clk), .RN(rst_n), .Q(
        conv_1[204]) );
  DFFRHQXL conv_1_reg_13__10_ ( .D(n16258), .CK(clk), .RN(rst_n), .Q(
        conv_1[205]) );
  DFFRHQXL conv_1_reg_13__11_ ( .D(n16257), .CK(clk), .RN(rst_n), .Q(
        conv_1[206]) );
  DFFRHQXL conv_1_reg_13__12_ ( .D(n16256), .CK(clk), .RN(rst_n), .Q(
        conv_1[207]) );
  DFFRHQXL conv_1_reg_13__13_ ( .D(n16255), .CK(clk), .RN(rst_n), .Q(
        conv_1[208]) );
  DFFRHQXL conv_1_reg_14__14_ ( .D(n16239), .CK(clk), .RN(rst_n), .Q(
        conv_1[224]) );
  DFFRHQXL conv_1_reg_14__0_ ( .D(n16253), .CK(clk), .RN(rst_n), .Q(
        conv_1[210]) );
  DFFRHQXL conv_1_reg_14__5_ ( .D(n16248), .CK(clk), .RN(rst_n), .Q(
        conv_1[215]) );
  DFFRHQXL conv_1_reg_14__6_ ( .D(n16247), .CK(clk), .RN(rst_n), .Q(
        conv_1[216]) );
  DFFRHQXL conv_1_reg_14__7_ ( .D(n16246), .CK(clk), .RN(rst_n), .Q(
        conv_1[217]) );
  DFFRHQXL conv_1_reg_14__8_ ( .D(n16245), .CK(clk), .RN(rst_n), .Q(
        conv_1[218]) );
  DFFRHQXL conv_1_reg_14__9_ ( .D(n16244), .CK(clk), .RN(rst_n), .Q(
        conv_1[219]) );
  DFFRHQXL conv_1_reg_14__10_ ( .D(n16243), .CK(clk), .RN(rst_n), .Q(
        conv_1[220]) );
  DFFRHQXL conv_1_reg_14__11_ ( .D(n16242), .CK(clk), .RN(rst_n), .Q(
        conv_1[221]) );
  DFFRHQXL conv_1_reg_14__12_ ( .D(n16241), .CK(clk), .RN(rst_n), .Q(
        conv_1[222]) );
  DFFRHQXL conv_1_reg_14__13_ ( .D(n16240), .CK(clk), .RN(rst_n), .Q(
        conv_1[223]) );
  DFFRHQXL conv_1_reg_15__14_ ( .D(n16224), .CK(clk), .RN(rst_n), .Q(
        conv_1[239]) );
  DFFRHQXL conv_1_reg_15__0_ ( .D(n16238), .CK(clk), .RN(rst_n), .Q(
        conv_1[225]) );
  DFFRHQXL conv_1_reg_15__5_ ( .D(n16233), .CK(clk), .RN(rst_n), .Q(
        conv_1[230]) );
  DFFRHQXL conv_1_reg_15__6_ ( .D(n16232), .CK(clk), .RN(rst_n), .Q(
        conv_1[231]) );
  DFFRHQXL conv_1_reg_15__7_ ( .D(n16231), .CK(clk), .RN(rst_n), .Q(
        conv_1[232]) );
  DFFRHQXL conv_1_reg_15__8_ ( .D(n16230), .CK(clk), .RN(rst_n), .Q(
        conv_1[233]) );
  DFFRHQXL conv_1_reg_15__9_ ( .D(n16229), .CK(clk), .RN(rst_n), .Q(
        conv_1[234]) );
  DFFRHQXL conv_1_reg_15__10_ ( .D(n16228), .CK(clk), .RN(rst_n), .Q(
        conv_1[235]) );
  DFFRHQXL conv_1_reg_15__11_ ( .D(n16227), .CK(clk), .RN(rst_n), .Q(
        conv_1[236]) );
  DFFRHQXL conv_1_reg_15__12_ ( .D(n16226), .CK(clk), .RN(rst_n), .Q(
        conv_1[237]) );
  DFFRHQXL conv_1_reg_15__13_ ( .D(n16225), .CK(clk), .RN(rst_n), .Q(
        conv_1[238]) );
  DFFRHQXL conv_1_reg_16__14_ ( .D(n16209), .CK(clk), .RN(rst_n), .Q(
        conv_1[254]) );
  DFFRHQXL conv_1_reg_16__0_ ( .D(n16223), .CK(clk), .RN(rst_n), .Q(
        conv_1[240]) );
  DFFRHQXL conv_1_reg_16__5_ ( .D(n16218), .CK(clk), .RN(rst_n), .Q(
        conv_1[245]) );
  DFFRHQXL conv_1_reg_16__6_ ( .D(n16217), .CK(clk), .RN(rst_n), .Q(
        conv_1[246]) );
  DFFRHQXL conv_1_reg_16__7_ ( .D(n16216), .CK(clk), .RN(rst_n), .Q(
        conv_1[247]) );
  DFFRHQXL conv_1_reg_16__8_ ( .D(n16215), .CK(clk), .RN(rst_n), .Q(
        conv_1[248]) );
  DFFRHQXL conv_1_reg_16__9_ ( .D(n16214), .CK(clk), .RN(rst_n), .Q(
        conv_1[249]) );
  DFFRHQXL conv_1_reg_16__10_ ( .D(n16213), .CK(clk), .RN(rst_n), .Q(
        conv_1[250]) );
  DFFRHQXL conv_1_reg_16__11_ ( .D(n16212), .CK(clk), .RN(rst_n), .Q(
        conv_1[251]) );
  DFFRHQXL conv_1_reg_16__12_ ( .D(n16211), .CK(clk), .RN(rst_n), .Q(
        conv_1[252]) );
  DFFRHQXL conv_1_reg_16__13_ ( .D(n16210), .CK(clk), .RN(rst_n), .Q(
        conv_1[253]) );
  DFFRHQXL conv_1_reg_17__14_ ( .D(n16194), .CK(clk), .RN(rst_n), .Q(
        conv_1[269]) );
  DFFRHQXL conv_1_reg_17__0_ ( .D(n16208), .CK(clk), .RN(rst_n), .Q(
        conv_1[255]) );
  DFFRHQXL conv_1_reg_17__5_ ( .D(n16203), .CK(clk), .RN(rst_n), .Q(
        conv_1[260]) );
  DFFRHQXL conv_1_reg_17__6_ ( .D(n16202), .CK(clk), .RN(rst_n), .Q(
        conv_1[261]) );
  DFFRHQXL conv_1_reg_17__7_ ( .D(n16201), .CK(clk), .RN(rst_n), .Q(
        conv_1[262]) );
  DFFRHQXL conv_1_reg_17__8_ ( .D(n16200), .CK(clk), .RN(rst_n), .Q(
        conv_1[263]) );
  DFFRHQXL conv_1_reg_17__9_ ( .D(n16199), .CK(clk), .RN(rst_n), .Q(
        conv_1[264]) );
  DFFRHQXL conv_1_reg_17__10_ ( .D(n16198), .CK(clk), .RN(rst_n), .Q(
        conv_1[265]) );
  DFFRHQXL conv_1_reg_17__11_ ( .D(n16197), .CK(clk), .RN(rst_n), .Q(
        conv_1[266]) );
  DFFRHQXL conv_1_reg_17__12_ ( .D(n16196), .CK(clk), .RN(rst_n), .Q(
        conv_1[267]) );
  DFFRHQXL conv_1_reg_17__13_ ( .D(n16195), .CK(clk), .RN(rst_n), .Q(
        conv_1[268]) );
  DFFRHQXL conv_1_reg_18__14_ ( .D(n16179), .CK(clk), .RN(rst_n), .Q(
        conv_1[284]) );
  DFFRHQXL conv_1_reg_18__0_ ( .D(n16193), .CK(clk), .RN(rst_n), .Q(
        conv_1[270]) );
  DFFRHQXL conv_1_reg_18__5_ ( .D(n16188), .CK(clk), .RN(rst_n), .Q(
        conv_1[275]) );
  DFFRHQXL conv_1_reg_18__6_ ( .D(n16187), .CK(clk), .RN(rst_n), .Q(
        conv_1[276]) );
  DFFRHQXL conv_1_reg_18__7_ ( .D(n16186), .CK(clk), .RN(rst_n), .Q(
        conv_1[277]) );
  DFFRHQXL conv_1_reg_18__8_ ( .D(n16185), .CK(clk), .RN(rst_n), .Q(
        conv_1[278]) );
  DFFRHQXL conv_1_reg_18__9_ ( .D(n16184), .CK(clk), .RN(rst_n), .Q(
        conv_1[279]) );
  DFFRHQXL conv_1_reg_18__10_ ( .D(n16183), .CK(clk), .RN(rst_n), .Q(
        conv_1[280]) );
  DFFRHQXL conv_1_reg_18__11_ ( .D(n16182), .CK(clk), .RN(rst_n), .Q(
        conv_1[281]) );
  DFFRHQXL conv_1_reg_18__12_ ( .D(n16181), .CK(clk), .RN(rst_n), .Q(
        conv_1[282]) );
  DFFRHQXL conv_1_reg_18__13_ ( .D(n16180), .CK(clk), .RN(rst_n), .Q(
        conv_1[283]) );
  DFFRHQXL conv_1_reg_19__14_ ( .D(n16164), .CK(clk), .RN(rst_n), .Q(
        conv_1[299]) );
  DFFRHQXL conv_1_reg_19__0_ ( .D(n16178), .CK(clk), .RN(rst_n), .Q(
        conv_1[285]) );
  DFFRHQXL conv_1_reg_19__5_ ( .D(n16173), .CK(clk), .RN(rst_n), .Q(
        conv_1[290]) );
  DFFRHQXL conv_1_reg_19__6_ ( .D(n16172), .CK(clk), .RN(rst_n), .Q(
        conv_1[291]) );
  DFFRHQXL conv_1_reg_19__7_ ( .D(n16171), .CK(clk), .RN(rst_n), .Q(
        conv_1[292]) );
  DFFRHQXL conv_1_reg_19__8_ ( .D(n16170), .CK(clk), .RN(rst_n), .Q(
        conv_1[293]) );
  DFFRHQXL conv_1_reg_19__9_ ( .D(n16169), .CK(clk), .RN(rst_n), .Q(
        conv_1[294]) );
  DFFRHQXL conv_1_reg_19__10_ ( .D(n16168), .CK(clk), .RN(rst_n), .Q(
        conv_1[295]) );
  DFFRHQXL conv_1_reg_19__11_ ( .D(n16167), .CK(clk), .RN(rst_n), .Q(
        conv_1[296]) );
  DFFRHQXL conv_1_reg_19__12_ ( .D(n16166), .CK(clk), .RN(rst_n), .Q(
        conv_1[297]) );
  DFFRHQXL conv_1_reg_19__13_ ( .D(n16165), .CK(clk), .RN(rst_n), .Q(
        conv_1[298]) );
  DFFRHQXL conv_1_reg_20__14_ ( .D(n16149), .CK(clk), .RN(rst_n), .Q(
        conv_1[314]) );
  DFFRHQXL conv_1_reg_20__0_ ( .D(n16163), .CK(clk), .RN(rst_n), .Q(
        conv_1[300]) );
  DFFRHQXL conv_1_reg_20__5_ ( .D(n16158), .CK(clk), .RN(rst_n), .Q(
        conv_1[305]) );
  DFFRHQXL conv_1_reg_20__6_ ( .D(n16157), .CK(clk), .RN(rst_n), .Q(
        conv_1[306]) );
  DFFRHQXL conv_1_reg_20__7_ ( .D(n16156), .CK(clk), .RN(rst_n), .Q(
        conv_1[307]) );
  DFFRHQXL conv_1_reg_20__8_ ( .D(n16155), .CK(clk), .RN(rst_n), .Q(
        conv_1[308]) );
  DFFRHQXL conv_1_reg_20__9_ ( .D(n16154), .CK(clk), .RN(rst_n), .Q(
        conv_1[309]) );
  DFFRHQXL conv_1_reg_20__10_ ( .D(n16153), .CK(clk), .RN(rst_n), .Q(
        conv_1[310]) );
  DFFRHQXL conv_1_reg_20__11_ ( .D(n16152), .CK(clk), .RN(rst_n), .Q(
        conv_1[311]) );
  DFFRHQXL conv_1_reg_20__12_ ( .D(n16151), .CK(clk), .RN(rst_n), .Q(
        conv_1[312]) );
  DFFRHQXL conv_1_reg_20__13_ ( .D(n16150), .CK(clk), .RN(rst_n), .Q(
        conv_1[313]) );
  DFFRHQXL conv_1_reg_21__14_ ( .D(n16134), .CK(clk), .RN(rst_n), .Q(
        conv_1[329]) );
  DFFRHQXL conv_1_reg_21__0_ ( .D(n16148), .CK(clk), .RN(rst_n), .Q(
        conv_1[315]) );
  DFFRHQXL conv_1_reg_21__5_ ( .D(n16143), .CK(clk), .RN(rst_n), .Q(
        conv_1[320]) );
  DFFRHQXL conv_1_reg_21__6_ ( .D(n16142), .CK(clk), .RN(rst_n), .Q(
        conv_1[321]) );
  DFFRHQXL conv_1_reg_21__7_ ( .D(n16141), .CK(clk), .RN(rst_n), .Q(
        conv_1[322]) );
  DFFRHQXL conv_1_reg_21__8_ ( .D(n16140), .CK(clk), .RN(rst_n), .Q(
        conv_1[323]) );
  DFFRHQXL conv_1_reg_21__9_ ( .D(n16139), .CK(clk), .RN(rst_n), .Q(
        conv_1[324]) );
  DFFRHQXL conv_1_reg_21__10_ ( .D(n16138), .CK(clk), .RN(rst_n), .Q(
        conv_1[325]) );
  DFFRHQXL conv_1_reg_21__11_ ( .D(n16137), .CK(clk), .RN(rst_n), .Q(
        conv_1[326]) );
  DFFRHQXL conv_1_reg_21__12_ ( .D(n16136), .CK(clk), .RN(rst_n), .Q(
        conv_1[327]) );
  DFFRHQXL conv_1_reg_21__13_ ( .D(n16135), .CK(clk), .RN(rst_n), .Q(
        conv_1[328]) );
  DFFRHQXL conv_1_reg_22__14_ ( .D(n16119), .CK(clk), .RN(rst_n), .Q(
        conv_1[344]) );
  DFFRHQXL conv_1_reg_22__0_ ( .D(n16133), .CK(clk), .RN(rst_n), .Q(
        conv_1[330]) );
  DFFRHQXL conv_1_reg_22__5_ ( .D(n16128), .CK(clk), .RN(rst_n), .Q(
        conv_1[335]) );
  DFFRHQXL conv_1_reg_22__6_ ( .D(n16127), .CK(clk), .RN(rst_n), .Q(
        conv_1[336]) );
  DFFRHQXL conv_1_reg_22__7_ ( .D(n16126), .CK(clk), .RN(rst_n), .Q(
        conv_1[337]) );
  DFFRHQXL conv_1_reg_22__8_ ( .D(n16125), .CK(clk), .RN(rst_n), .Q(
        conv_1[338]) );
  DFFRHQXL conv_1_reg_22__9_ ( .D(n16124), .CK(clk), .RN(rst_n), .Q(
        conv_1[339]) );
  DFFRHQXL conv_1_reg_22__10_ ( .D(n16123), .CK(clk), .RN(rst_n), .Q(
        conv_1[340]) );
  DFFRHQXL conv_1_reg_22__11_ ( .D(n16122), .CK(clk), .RN(rst_n), .Q(
        conv_1[341]) );
  DFFRHQXL conv_1_reg_22__12_ ( .D(n16121), .CK(clk), .RN(rst_n), .Q(
        conv_1[342]) );
  DFFRHQXL conv_1_reg_22__13_ ( .D(n16120), .CK(clk), .RN(rst_n), .Q(
        conv_1[343]) );
  DFFRHQXL conv_1_reg_23__14_ ( .D(n16104), .CK(clk), .RN(rst_n), .Q(
        conv_1[359]) );
  DFFRHQXL conv_1_reg_23__0_ ( .D(n16118), .CK(clk), .RN(rst_n), .Q(
        conv_1[345]) );
  DFFRHQXL conv_1_reg_23__5_ ( .D(n16113), .CK(clk), .RN(rst_n), .Q(
        conv_1[350]) );
  DFFRHQXL conv_1_reg_23__6_ ( .D(n16112), .CK(clk), .RN(rst_n), .Q(
        conv_1[351]) );
  DFFRHQXL conv_1_reg_23__7_ ( .D(n16111), .CK(clk), .RN(rst_n), .Q(
        conv_1[352]) );
  DFFRHQXL conv_1_reg_23__8_ ( .D(n16110), .CK(clk), .RN(rst_n), .Q(
        conv_1[353]) );
  DFFRHQXL conv_1_reg_23__9_ ( .D(n16109), .CK(clk), .RN(rst_n), .Q(
        conv_1[354]) );
  DFFRHQXL conv_1_reg_23__10_ ( .D(n16108), .CK(clk), .RN(rst_n), .Q(
        conv_1[355]) );
  DFFRHQXL conv_1_reg_23__11_ ( .D(n16107), .CK(clk), .RN(rst_n), .Q(
        conv_1[356]) );
  DFFRHQXL conv_1_reg_23__12_ ( .D(n16106), .CK(clk), .RN(rst_n), .Q(
        conv_1[357]) );
  DFFRHQXL conv_1_reg_23__13_ ( .D(n16105), .CK(clk), .RN(rst_n), .Q(
        conv_1[358]) );
  DFFRHQXL conv_1_reg_24__14_ ( .D(n16089), .CK(clk), .RN(rst_n), .Q(
        conv_1[374]) );
  DFFRHQXL conv_1_reg_24__0_ ( .D(n16103), .CK(clk), .RN(rst_n), .Q(
        conv_1[360]) );
  DFFRHQXL conv_1_reg_24__5_ ( .D(n16098), .CK(clk), .RN(rst_n), .Q(
        conv_1[365]) );
  DFFRHQXL conv_1_reg_24__6_ ( .D(n16097), .CK(clk), .RN(rst_n), .Q(
        conv_1[366]) );
  DFFRHQXL conv_1_reg_24__7_ ( .D(n16096), .CK(clk), .RN(rst_n), .Q(
        conv_1[367]) );
  DFFRHQXL conv_1_reg_24__8_ ( .D(n16095), .CK(clk), .RN(rst_n), .Q(
        conv_1[368]) );
  DFFRHQXL conv_1_reg_24__9_ ( .D(n16094), .CK(clk), .RN(rst_n), .Q(
        conv_1[369]) );
  DFFRHQXL conv_1_reg_24__10_ ( .D(n16093), .CK(clk), .RN(rst_n), .Q(
        conv_1[370]) );
  DFFRHQXL conv_1_reg_24__11_ ( .D(n16092), .CK(clk), .RN(rst_n), .Q(
        conv_1[371]) );
  DFFRHQXL conv_1_reg_24__12_ ( .D(n16091), .CK(clk), .RN(rst_n), .Q(
        conv_1[372]) );
  DFFRHQXL conv_1_reg_24__13_ ( .D(n16090), .CK(clk), .RN(rst_n), .Q(
        conv_1[373]) );
  DFFRHQXL conv_1_reg_25__14_ ( .D(n16074), .CK(clk), .RN(rst_n), .Q(
        conv_1[389]) );
  DFFRHQXL conv_1_reg_25__0_ ( .D(n16088), .CK(clk), .RN(rst_n), .Q(
        conv_1[375]) );
  DFFRHQXL conv_1_reg_25__5_ ( .D(n16083), .CK(clk), .RN(rst_n), .Q(
        conv_1[380]) );
  DFFRHQXL conv_1_reg_25__6_ ( .D(n16082), .CK(clk), .RN(rst_n), .Q(
        conv_1[381]) );
  DFFRHQXL conv_1_reg_25__7_ ( .D(n16081), .CK(clk), .RN(rst_n), .Q(
        conv_1[382]) );
  DFFRHQXL conv_1_reg_25__8_ ( .D(n16080), .CK(clk), .RN(rst_n), .Q(
        conv_1[383]) );
  DFFRHQXL conv_1_reg_25__9_ ( .D(n16079), .CK(clk), .RN(rst_n), .Q(
        conv_1[384]) );
  DFFRHQXL conv_1_reg_25__10_ ( .D(n16078), .CK(clk), .RN(rst_n), .Q(
        conv_1[385]) );
  DFFRHQXL conv_1_reg_25__11_ ( .D(n16077), .CK(clk), .RN(rst_n), .Q(
        conv_1[386]) );
  DFFRHQXL conv_1_reg_25__12_ ( .D(n16076), .CK(clk), .RN(rst_n), .Q(
        conv_1[387]) );
  DFFRHQXL conv_1_reg_25__13_ ( .D(n16075), .CK(clk), .RN(rst_n), .Q(
        conv_1[388]) );
  DFFRHQXL conv_1_reg_26__14_ ( .D(n16059), .CK(clk), .RN(rst_n), .Q(
        conv_1[404]) );
  DFFRHQXL conv_1_reg_26__0_ ( .D(n16073), .CK(clk), .RN(rst_n), .Q(
        conv_1[390]) );
  DFFRHQXL conv_1_reg_26__5_ ( .D(n16068), .CK(clk), .RN(rst_n), .Q(
        conv_1[395]) );
  DFFRHQXL conv_1_reg_26__6_ ( .D(n16067), .CK(clk), .RN(rst_n), .Q(
        conv_1[396]) );
  DFFRHQXL conv_1_reg_26__7_ ( .D(n16066), .CK(clk), .RN(rst_n), .Q(
        conv_1[397]) );
  DFFRHQXL conv_1_reg_26__8_ ( .D(n16065), .CK(clk), .RN(rst_n), .Q(
        conv_1[398]) );
  DFFRHQXL conv_1_reg_26__9_ ( .D(n16064), .CK(clk), .RN(rst_n), .Q(
        conv_1[399]) );
  DFFRHQXL conv_1_reg_26__10_ ( .D(n16063), .CK(clk), .RN(rst_n), .Q(
        conv_1[400]) );
  DFFRHQXL conv_1_reg_26__11_ ( .D(n16062), .CK(clk), .RN(rst_n), .Q(
        conv_1[401]) );
  DFFRHQXL conv_1_reg_26__12_ ( .D(n16061), .CK(clk), .RN(rst_n), .Q(
        conv_1[402]) );
  DFFRHQXL conv_1_reg_26__13_ ( .D(n16060), .CK(clk), .RN(rst_n), .Q(
        conv_1[403]) );
  DFFRHQXL conv_1_reg_27__14_ ( .D(n16044), .CK(clk), .RN(rst_n), .Q(
        conv_1[419]) );
  DFFRHQXL conv_1_reg_27__0_ ( .D(n16058), .CK(clk), .RN(rst_n), .Q(
        conv_1[405]) );
  DFFRHQXL conv_1_reg_27__5_ ( .D(n16053), .CK(clk), .RN(rst_n), .Q(
        conv_1[410]) );
  DFFRHQXL conv_1_reg_27__6_ ( .D(n16052), .CK(clk), .RN(rst_n), .Q(
        conv_1[411]) );
  DFFRHQXL conv_1_reg_27__7_ ( .D(n16051), .CK(clk), .RN(rst_n), .Q(
        conv_1[412]) );
  DFFRHQXL conv_1_reg_27__8_ ( .D(n16050), .CK(clk), .RN(rst_n), .Q(
        conv_1[413]) );
  DFFRHQXL conv_1_reg_27__9_ ( .D(n16049), .CK(clk), .RN(rst_n), .Q(
        conv_1[414]) );
  DFFRHQXL conv_1_reg_27__10_ ( .D(n16048), .CK(clk), .RN(rst_n), .Q(
        conv_1[415]) );
  DFFRHQXL conv_1_reg_27__11_ ( .D(n16047), .CK(clk), .RN(rst_n), .Q(
        conv_1[416]) );
  DFFRHQXL conv_1_reg_27__12_ ( .D(n16046), .CK(clk), .RN(rst_n), .Q(
        conv_1[417]) );
  DFFRHQXL conv_1_reg_27__13_ ( .D(n16045), .CK(clk), .RN(rst_n), .Q(
        conv_1[418]) );
  DFFRHQXL conv_1_reg_28__14_ ( .D(n16029), .CK(clk), .RN(rst_n), .Q(
        conv_1[434]) );
  DFFRHQXL conv_1_reg_28__0_ ( .D(n16043), .CK(clk), .RN(rst_n), .Q(
        conv_1[420]) );
  DFFRHQXL conv_1_reg_28__5_ ( .D(n16038), .CK(clk), .RN(rst_n), .Q(
        conv_1[425]) );
  DFFRHQXL conv_1_reg_28__6_ ( .D(n16037), .CK(clk), .RN(rst_n), .Q(
        conv_1[426]) );
  DFFRHQXL conv_1_reg_28__7_ ( .D(n16036), .CK(clk), .RN(rst_n), .Q(
        conv_1[427]) );
  DFFRHQXL conv_1_reg_28__8_ ( .D(n16035), .CK(clk), .RN(rst_n), .Q(
        conv_1[428]) );
  DFFRHQXL conv_1_reg_28__9_ ( .D(n16034), .CK(clk), .RN(rst_n), .Q(
        conv_1[429]) );
  DFFRHQXL conv_1_reg_28__10_ ( .D(n16033), .CK(clk), .RN(rst_n), .Q(
        conv_1[430]) );
  DFFRHQXL conv_1_reg_28__11_ ( .D(n16032), .CK(clk), .RN(rst_n), .Q(
        conv_1[431]) );
  DFFRHQXL conv_1_reg_28__12_ ( .D(n16031), .CK(clk), .RN(rst_n), .Q(
        conv_1[432]) );
  DFFRHQXL conv_1_reg_28__13_ ( .D(n16030), .CK(clk), .RN(rst_n), .Q(
        conv_1[433]) );
  DFFRHQXL conv_1_reg_29__14_ ( .D(n16014), .CK(clk), .RN(rst_n), .Q(
        conv_1[449]) );
  DFFRHQXL conv_1_reg_29__0_ ( .D(n16028), .CK(clk), .RN(rst_n), .Q(
        conv_1[435]) );
  DFFRHQXL conv_1_reg_29__5_ ( .D(n16023), .CK(clk), .RN(rst_n), .Q(
        conv_1[440]) );
  DFFRHQXL conv_1_reg_29__6_ ( .D(n16022), .CK(clk), .RN(rst_n), .Q(
        conv_1[441]) );
  DFFRHQXL conv_1_reg_29__7_ ( .D(n16021), .CK(clk), .RN(rst_n), .Q(
        conv_1[442]) );
  DFFRHQXL conv_1_reg_29__8_ ( .D(n16020), .CK(clk), .RN(rst_n), .Q(
        conv_1[443]) );
  DFFRHQXL conv_1_reg_29__9_ ( .D(n16019), .CK(clk), .RN(rst_n), .Q(
        conv_1[444]) );
  DFFRHQXL conv_1_reg_29__10_ ( .D(n16018), .CK(clk), .RN(rst_n), .Q(
        conv_1[445]) );
  DFFRHQXL conv_1_reg_29__11_ ( .D(n16017), .CK(clk), .RN(rst_n), .Q(
        conv_1[446]) );
  DFFRHQXL conv_1_reg_29__12_ ( .D(n16016), .CK(clk), .RN(rst_n), .Q(
        conv_1[447]) );
  DFFRHQXL conv_1_reg_29__13_ ( .D(n16015), .CK(clk), .RN(rst_n), .Q(
        conv_1[448]) );
  DFFRHQXL conv_1_reg_30__14_ ( .D(n15999), .CK(clk), .RN(rst_n), .Q(
        conv_1[464]) );
  DFFRHQXL conv_1_reg_30__0_ ( .D(n16013), .CK(clk), .RN(rst_n), .Q(
        conv_1[450]) );
  DFFRHQXL conv_1_reg_30__5_ ( .D(n16008), .CK(clk), .RN(rst_n), .Q(
        conv_1[455]) );
  DFFRHQXL conv_1_reg_30__6_ ( .D(n16007), .CK(clk), .RN(rst_n), .Q(
        conv_1[456]) );
  DFFRHQXL conv_1_reg_30__7_ ( .D(n16006), .CK(clk), .RN(rst_n), .Q(
        conv_1[457]) );
  DFFRHQXL conv_1_reg_30__8_ ( .D(n16005), .CK(clk), .RN(rst_n), .Q(
        conv_1[458]) );
  DFFRHQXL conv_1_reg_30__9_ ( .D(n16004), .CK(clk), .RN(rst_n), .Q(
        conv_1[459]) );
  DFFRHQXL conv_1_reg_30__10_ ( .D(n16003), .CK(clk), .RN(rst_n), .Q(
        conv_1[460]) );
  DFFRHQXL conv_1_reg_30__11_ ( .D(n16002), .CK(clk), .RN(rst_n), .Q(
        conv_1[461]) );
  DFFRHQXL conv_1_reg_30__12_ ( .D(n16001), .CK(clk), .RN(rst_n), .Q(
        conv_1[462]) );
  DFFRHQXL conv_1_reg_30__13_ ( .D(n16000), .CK(clk), .RN(rst_n), .Q(
        conv_1[463]) );
  DFFRHQXL conv_1_reg_31__14_ ( .D(n15984), .CK(clk), .RN(rst_n), .Q(
        conv_1[479]) );
  DFFRHQXL conv_1_reg_31__0_ ( .D(n15998), .CK(clk), .RN(rst_n), .Q(
        conv_1[465]) );
  DFFRHQXL conv_1_reg_31__5_ ( .D(n15993), .CK(clk), .RN(rst_n), .Q(
        conv_1[470]) );
  DFFRHQXL conv_1_reg_31__6_ ( .D(n15992), .CK(clk), .RN(rst_n), .Q(
        conv_1[471]) );
  DFFRHQXL conv_1_reg_31__7_ ( .D(n15991), .CK(clk), .RN(rst_n), .Q(
        conv_1[472]) );
  DFFRHQXL conv_1_reg_31__8_ ( .D(n15990), .CK(clk), .RN(rst_n), .Q(
        conv_1[473]) );
  DFFRHQXL conv_1_reg_31__9_ ( .D(n15989), .CK(clk), .RN(rst_n), .Q(
        conv_1[474]) );
  DFFRHQXL conv_1_reg_31__10_ ( .D(n15988), .CK(clk), .RN(rst_n), .Q(
        conv_1[475]) );
  DFFRHQXL conv_1_reg_31__11_ ( .D(n15987), .CK(clk), .RN(rst_n), .Q(
        conv_1[476]) );
  DFFRHQXL conv_1_reg_31__12_ ( .D(n15986), .CK(clk), .RN(rst_n), .Q(
        conv_1[477]) );
  DFFRHQXL conv_1_reg_31__13_ ( .D(n15985), .CK(clk), .RN(rst_n), .Q(
        conv_1[478]) );
  DFFRHQXL conv_1_reg_32__14_ ( .D(n15969), .CK(clk), .RN(rst_n), .Q(
        conv_1[494]) );
  DFFRHQXL conv_1_reg_32__0_ ( .D(n15983), .CK(clk), .RN(rst_n), .Q(
        conv_1[480]) );
  DFFRHQXL conv_1_reg_32__5_ ( .D(n15978), .CK(clk), .RN(rst_n), .Q(
        conv_1[485]) );
  DFFRHQXL conv_1_reg_32__6_ ( .D(n15977), .CK(clk), .RN(rst_n), .Q(
        conv_1[486]) );
  DFFRHQXL conv_1_reg_32__7_ ( .D(n15976), .CK(clk), .RN(rst_n), .Q(
        conv_1[487]) );
  DFFRHQXL conv_1_reg_32__8_ ( .D(n15975), .CK(clk), .RN(rst_n), .Q(
        conv_1[488]) );
  DFFRHQXL conv_1_reg_32__9_ ( .D(n15974), .CK(clk), .RN(rst_n), .Q(
        conv_1[489]) );
  DFFRHQXL conv_1_reg_32__10_ ( .D(n15973), .CK(clk), .RN(rst_n), .Q(
        conv_1[490]) );
  DFFRHQXL conv_1_reg_32__11_ ( .D(n15972), .CK(clk), .RN(rst_n), .Q(
        conv_1[491]) );
  DFFRHQXL conv_1_reg_32__12_ ( .D(n15971), .CK(clk), .RN(rst_n), .Q(
        conv_1[492]) );
  DFFRHQXL conv_1_reg_32__13_ ( .D(n15970), .CK(clk), .RN(rst_n), .Q(
        conv_1[493]) );
  DFFRHQXL conv_1_reg_33__14_ ( .D(n15954), .CK(clk), .RN(rst_n), .Q(
        conv_1[509]) );
  DFFRHQXL conv_1_reg_33__0_ ( .D(n15968), .CK(clk), .RN(rst_n), .Q(
        conv_1[495]) );
  DFFRHQXL conv_1_reg_33__5_ ( .D(n15963), .CK(clk), .RN(rst_n), .Q(
        conv_1[500]) );
  DFFRHQXL conv_1_reg_33__6_ ( .D(n15962), .CK(clk), .RN(rst_n), .Q(
        conv_1[501]) );
  DFFRHQXL conv_1_reg_33__7_ ( .D(n15961), .CK(clk), .RN(rst_n), .Q(
        conv_1[502]) );
  DFFRHQXL conv_1_reg_33__8_ ( .D(n15960), .CK(clk), .RN(rst_n), .Q(
        conv_1[503]) );
  DFFRHQXL conv_1_reg_33__9_ ( .D(n15959), .CK(clk), .RN(rst_n), .Q(
        conv_1[504]) );
  DFFRHQXL conv_1_reg_33__10_ ( .D(n15958), .CK(clk), .RN(rst_n), .Q(
        conv_1[505]) );
  DFFRHQXL conv_1_reg_33__11_ ( .D(n15957), .CK(clk), .RN(rst_n), .Q(
        conv_1[506]) );
  DFFRHQXL conv_1_reg_33__12_ ( .D(n15956), .CK(clk), .RN(rst_n), .Q(
        conv_1[507]) );
  DFFRHQXL conv_1_reg_33__13_ ( .D(n15955), .CK(clk), .RN(rst_n), .Q(
        conv_1[508]) );
  DFFRHQXL conv_1_reg_34__14_ ( .D(n15939), .CK(clk), .RN(rst_n), .Q(
        conv_1[524]) );
  DFFRHQXL conv_1_reg_34__0_ ( .D(n15953), .CK(clk), .RN(rst_n), .Q(
        conv_1[510]) );
  DFFRHQXL conv_1_reg_34__5_ ( .D(n15948), .CK(clk), .RN(rst_n), .Q(
        conv_1[515]) );
  DFFRHQXL conv_1_reg_34__6_ ( .D(n15947), .CK(clk), .RN(rst_n), .Q(
        conv_1[516]) );
  DFFRHQXL conv_1_reg_34__7_ ( .D(n15946), .CK(clk), .RN(rst_n), .Q(
        conv_1[517]) );
  DFFRHQXL conv_1_reg_34__8_ ( .D(n15945), .CK(clk), .RN(rst_n), .Q(
        conv_1[518]) );
  DFFRHQXL conv_1_reg_34__9_ ( .D(n15944), .CK(clk), .RN(rst_n), .Q(
        conv_1[519]) );
  DFFRHQXL conv_1_reg_34__10_ ( .D(n15943), .CK(clk), .RN(rst_n), .Q(
        conv_1[520]) );
  DFFRHQXL conv_1_reg_34__11_ ( .D(n15942), .CK(clk), .RN(rst_n), .Q(
        conv_1[521]) );
  DFFRHQXL conv_1_reg_34__12_ ( .D(n15941), .CK(clk), .RN(rst_n), .Q(
        conv_1[522]) );
  DFFRHQXL conv_1_reg_34__13_ ( .D(n15940), .CK(clk), .RN(rst_n), .Q(
        conv_1[523]) );
  DFFRHQXL conv_1_reg_35__14_ ( .D(n15924), .CK(clk), .RN(rst_n), .Q(
        conv_1[539]) );
  DFFRHQXL conv_1_reg_35__0_ ( .D(n15938), .CK(clk), .RN(rst_n), .Q(
        conv_1[525]) );
  DFFRHQXL pool_reg_6__0_ ( .D(N29246), .CK(clk), .RN(rst_n), .Q(pool[30]) );
  DFFRHQXL pool_reg_8__0_ ( .D(N29256), .CK(clk), .RN(rst_n), .Q(pool[40]) );
  DFFRHQXL pool_reg_3__0_ ( .D(N29231), .CK(clk), .RN(rst_n), .Q(pool[15]) );
  DFFRHQXL pool_reg_2__0_ ( .D(N29226), .CK(clk), .RN(rst_n), .Q(pool[10]) );
  DFFRHQXL pool_reg_5__0_ ( .D(N29241), .CK(clk), .RN(rst_n), .Q(pool[25]) );
  DFFRHQXL pool_reg_0__0_ ( .D(N29216), .CK(clk), .RN(rst_n), .Q(pool[0]) );
  DFFRHQXL pool_reg_1__0_ ( .D(N29221), .CK(clk), .RN(rst_n), .Q(pool[5]) );
  DFFRHQXL pool_reg_7__0_ ( .D(N29251), .CK(clk), .RN(rst_n), .Q(pool[35]) );
  DFFRHQXL pool_reg_4__0_ ( .D(N29236), .CK(clk), .RN(rst_n), .Q(pool[20]) );
  DFFRHQXL conv_1_reg_35__5_ ( .D(n15933), .CK(clk), .RN(rst_n), .Q(
        conv_1[530]) );
  DFFRHQXL conv_1_reg_35__6_ ( .D(n15932), .CK(clk), .RN(rst_n), .Q(
        conv_1[531]) );
  DFFRHQXL conv_1_reg_35__7_ ( .D(n15931), .CK(clk), .RN(rst_n), .Q(
        conv_1[532]) );
  DFFRHQXL conv_1_reg_35__8_ ( .D(n15930), .CK(clk), .RN(rst_n), .Q(
        conv_1[533]) );
  DFFRHQXL conv_1_reg_35__9_ ( .D(n15929), .CK(clk), .RN(rst_n), .Q(
        conv_1[534]) );
  DFFRHQXL conv_1_reg_35__10_ ( .D(n15928), .CK(clk), .RN(rst_n), .Q(
        conv_1[535]) );
  DFFRHQXL conv_1_reg_35__11_ ( .D(n15927), .CK(clk), .RN(rst_n), .Q(
        conv_1[536]) );
  DFFRHQXL conv_1_reg_35__12_ ( .D(n15926), .CK(clk), .RN(rst_n), .Q(
        conv_1[537]) );
  DFFRHQXL conv_1_reg_35__13_ ( .D(n15925), .CK(clk), .RN(rst_n), .Q(
        conv_1[538]) );
  DFFRHQXL filter_3_bias_reg_4_ ( .D(n14729), .CK(clk), .RN(rst_n), .Q(
        filter_3_bias[4]) );
  DFFRHQXL conv_3_reg_0__4_ ( .D(n15779), .CK(clk), .RN(rst_n), .Q(conv_3[4])
         );
  DFFRHQXL conv_3_reg_1__4_ ( .D(n15778), .CK(clk), .RN(rst_n), .Q(conv_3[19])
         );
  DFFRHQXL conv_3_reg_2__4_ ( .D(n15777), .CK(clk), .RN(rst_n), .Q(conv_3[34])
         );
  DFFRHQXL conv_3_reg_3__4_ ( .D(n15776), .CK(clk), .RN(rst_n), .Q(conv_3[49])
         );
  DFFRHQXL conv_3_reg_4__4_ ( .D(n15775), .CK(clk), .RN(rst_n), .Q(conv_3[64])
         );
  DFFRHQXL conv_3_reg_5__4_ ( .D(n15774), .CK(clk), .RN(rst_n), .Q(conv_3[79])
         );
  DFFRHQXL conv_3_reg_6__4_ ( .D(n15773), .CK(clk), .RN(rst_n), .Q(conv_3[94])
         );
  DFFRHQXL conv_3_reg_7__4_ ( .D(n15772), .CK(clk), .RN(rst_n), .Q(conv_3[109]) );
  DFFRHQXL conv_3_reg_8__4_ ( .D(n15771), .CK(clk), .RN(rst_n), .Q(conv_3[124]) );
  DFFRHQXL conv_3_reg_9__4_ ( .D(n15770), .CK(clk), .RN(rst_n), .Q(conv_3[139]) );
  DFFRHQXL conv_3_reg_10__4_ ( .D(n15769), .CK(clk), .RN(rst_n), .Q(
        conv_3[154]) );
  DFFRHQXL conv_3_reg_11__4_ ( .D(n15768), .CK(clk), .RN(rst_n), .Q(
        conv_3[169]) );
  DFFRHQXL conv_3_reg_12__4_ ( .D(n15767), .CK(clk), .RN(rst_n), .Q(
        conv_3[184]) );
  DFFRHQXL conv_3_reg_13__4_ ( .D(n15766), .CK(clk), .RN(rst_n), .Q(
        conv_3[199]) );
  DFFRHQXL conv_3_reg_14__4_ ( .D(n15765), .CK(clk), .RN(rst_n), .Q(
        conv_3[214]) );
  DFFRHQXL conv_3_reg_15__4_ ( .D(n15764), .CK(clk), .RN(rst_n), .Q(
        conv_3[229]) );
  DFFRHQXL conv_3_reg_16__4_ ( .D(n15763), .CK(clk), .RN(rst_n), .Q(
        conv_3[244]) );
  DFFRHQXL conv_3_reg_17__4_ ( .D(n15762), .CK(clk), .RN(rst_n), .Q(
        conv_3[259]) );
  DFFRHQXL conv_3_reg_18__4_ ( .D(n15761), .CK(clk), .RN(rst_n), .Q(
        conv_3[274]) );
  DFFRHQXL conv_3_reg_19__4_ ( .D(n15760), .CK(clk), .RN(rst_n), .Q(
        conv_3[289]) );
  DFFRHQXL conv_3_reg_20__4_ ( .D(n15759), .CK(clk), .RN(rst_n), .Q(
        conv_3[304]) );
  DFFRHQXL conv_3_reg_21__4_ ( .D(n15758), .CK(clk), .RN(rst_n), .Q(
        conv_3[319]) );
  DFFRHQXL conv_3_reg_22__4_ ( .D(n15757), .CK(clk), .RN(rst_n), .Q(
        conv_3[334]) );
  DFFRHQXL conv_3_reg_23__4_ ( .D(n15756), .CK(clk), .RN(rst_n), .Q(
        conv_3[349]) );
  DFFRHQXL conv_3_reg_24__4_ ( .D(n15755), .CK(clk), .RN(rst_n), .Q(
        conv_3[364]) );
  DFFRHQXL conv_3_reg_25__4_ ( .D(n15754), .CK(clk), .RN(rst_n), .Q(
        conv_3[379]) );
  DFFRHQXL conv_3_reg_26__4_ ( .D(n15753), .CK(clk), .RN(rst_n), .Q(
        conv_3[394]) );
  DFFRHQXL conv_3_reg_27__4_ ( .D(n15752), .CK(clk), .RN(rst_n), .Q(
        conv_3[409]) );
  DFFRHQXL conv_3_reg_28__4_ ( .D(n15751), .CK(clk), .RN(rst_n), .Q(
        conv_3[424]) );
  DFFRHQXL conv_3_reg_29__4_ ( .D(n15750), .CK(clk), .RN(rst_n), .Q(
        conv_3[439]) );
  DFFRHQXL conv_3_reg_30__4_ ( .D(n15749), .CK(clk), .RN(rst_n), .Q(
        conv_3[454]) );
  DFFRHQXL conv_3_reg_31__4_ ( .D(n15748), .CK(clk), .RN(rst_n), .Q(
        conv_3[469]) );
  DFFRHQXL conv_3_reg_32__4_ ( .D(n15747), .CK(clk), .RN(rst_n), .Q(
        conv_3[484]) );
  DFFRHQXL conv_3_reg_33__4_ ( .D(n15746), .CK(clk), .RN(rst_n), .Q(
        conv_3[499]) );
  DFFRHQXL conv_3_reg_34__4_ ( .D(n15745), .CK(clk), .RN(rst_n), .Q(
        conv_3[514]) );
  DFFRHQXL conv_3_reg_35__4_ ( .D(n15744), .CK(clk), .RN(rst_n), .Q(
        conv_3[529]) );
  DFFRHQXL pool_reg_24__4_ ( .D(N29340), .CK(clk), .RN(rst_n), .Q(pool[124])
         );
  DFFRHQXL pool_reg_26__4_ ( .D(N29350), .CK(clk), .RN(rst_n), .Q(pool[134])
         );
  DFFRHQXL pool_reg_21__4_ ( .D(N29325), .CK(clk), .RN(rst_n), .Q(pool[109])
         );
  DFFRHQXL pool_reg_20__4_ ( .D(N29320), .CK(clk), .RN(rst_n), .Q(pool[104])
         );
  DFFRHQXL pool_reg_23__4_ ( .D(N29335), .CK(clk), .RN(rst_n), .Q(pool[119])
         );
  DFFRHQXL pool_reg_18__4_ ( .D(N29310), .CK(clk), .RN(rst_n), .Q(pool[94]) );
  DFFRHQXL pool_reg_19__4_ ( .D(N29315), .CK(clk), .RN(rst_n), .Q(pool[99]) );
  DFFRHQXL pool_reg_25__4_ ( .D(N29345), .CK(clk), .RN(rst_n), .Q(pool[129])
         );
  DFFRHQXL pool_reg_22__4_ ( .D(N29330), .CK(clk), .RN(rst_n), .Q(pool[114])
         );
  DFFRHQXL filter_2_bias_reg_4_ ( .D(n14728), .CK(clk), .RN(rst_n), .Q(
        filter_2_bias[4]) );
  DFFRHQXL conv_2_reg_0__4_ ( .D(n15239), .CK(clk), .RN(rst_n), .Q(conv_2[4])
         );
  DFFRHQXL conv_2_reg_1__4_ ( .D(n15238), .CK(clk), .RN(rst_n), .Q(conv_2[19])
         );
  DFFRHQXL conv_2_reg_2__4_ ( .D(n15237), .CK(clk), .RN(rst_n), .Q(conv_2[34])
         );
  DFFRHQXL conv_2_reg_3__4_ ( .D(n15236), .CK(clk), .RN(rst_n), .Q(conv_2[49])
         );
  DFFRHQXL conv_2_reg_4__4_ ( .D(n15235), .CK(clk), .RN(rst_n), .Q(conv_2[64])
         );
  DFFRHQXL conv_2_reg_5__4_ ( .D(n15234), .CK(clk), .RN(rst_n), .Q(conv_2[79])
         );
  DFFRHQXL conv_2_reg_6__4_ ( .D(n15233), .CK(clk), .RN(rst_n), .Q(conv_2[94])
         );
  DFFRHQXL conv_2_reg_7__4_ ( .D(n15232), .CK(clk), .RN(rst_n), .Q(conv_2[109]) );
  DFFRHQXL conv_2_reg_8__4_ ( .D(n15231), .CK(clk), .RN(rst_n), .Q(conv_2[124]) );
  DFFRHQXL conv_2_reg_9__4_ ( .D(n15230), .CK(clk), .RN(rst_n), .Q(conv_2[139]) );
  DFFRHQXL conv_2_reg_10__4_ ( .D(n15229), .CK(clk), .RN(rst_n), .Q(
        conv_2[154]) );
  DFFRHQXL conv_2_reg_11__4_ ( .D(n15228), .CK(clk), .RN(rst_n), .Q(
        conv_2[169]) );
  DFFRHQXL conv_2_reg_12__4_ ( .D(n15227), .CK(clk), .RN(rst_n), .Q(
        conv_2[184]) );
  DFFRHQXL conv_2_reg_13__4_ ( .D(n15226), .CK(clk), .RN(rst_n), .Q(
        conv_2[199]) );
  DFFRHQXL conv_2_reg_14__4_ ( .D(n15225), .CK(clk), .RN(rst_n), .Q(
        conv_2[214]) );
  DFFRHQXL conv_2_reg_15__4_ ( .D(n15224), .CK(clk), .RN(rst_n), .Q(
        conv_2[229]) );
  DFFRHQXL conv_2_reg_16__4_ ( .D(n15223), .CK(clk), .RN(rst_n), .Q(
        conv_2[244]) );
  DFFRHQXL conv_2_reg_17__4_ ( .D(n15222), .CK(clk), .RN(rst_n), .Q(
        conv_2[259]) );
  DFFRHQXL conv_2_reg_18__4_ ( .D(n15221), .CK(clk), .RN(rst_n), .Q(
        conv_2[274]) );
  DFFRHQXL conv_2_reg_19__4_ ( .D(n15220), .CK(clk), .RN(rst_n), .Q(
        conv_2[289]) );
  DFFRHQXL conv_2_reg_20__4_ ( .D(n15219), .CK(clk), .RN(rst_n), .Q(
        conv_2[304]) );
  DFFRHQXL conv_2_reg_21__4_ ( .D(n15218), .CK(clk), .RN(rst_n), .Q(
        conv_2[319]) );
  DFFRHQXL conv_2_reg_22__4_ ( .D(n15217), .CK(clk), .RN(rst_n), .Q(
        conv_2[334]) );
  DFFRHQXL conv_2_reg_23__4_ ( .D(n15216), .CK(clk), .RN(rst_n), .Q(
        conv_2[349]) );
  DFFRHQXL conv_2_reg_24__4_ ( .D(n15215), .CK(clk), .RN(rst_n), .Q(
        conv_2[364]) );
  DFFRHQXL conv_2_reg_25__4_ ( .D(n15214), .CK(clk), .RN(rst_n), .Q(
        conv_2[379]) );
  DFFRHQXL conv_2_reg_26__4_ ( .D(n15213), .CK(clk), .RN(rst_n), .Q(
        conv_2[394]) );
  DFFRHQXL conv_2_reg_27__4_ ( .D(n15212), .CK(clk), .RN(rst_n), .Q(
        conv_2[409]) );
  DFFRHQXL conv_2_reg_28__4_ ( .D(n15211), .CK(clk), .RN(rst_n), .Q(
        conv_2[424]) );
  DFFRHQXL conv_2_reg_29__4_ ( .D(n15210), .CK(clk), .RN(rst_n), .Q(
        conv_2[439]) );
  DFFRHQXL conv_2_reg_30__4_ ( .D(n15209), .CK(clk), .RN(rst_n), .Q(
        conv_2[454]) );
  DFFRHQXL conv_2_reg_31__4_ ( .D(n15208), .CK(clk), .RN(rst_n), .Q(
        conv_2[469]) );
  DFFRHQXL conv_2_reg_32__4_ ( .D(n15207), .CK(clk), .RN(rst_n), .Q(
        conv_2[484]) );
  DFFRHQXL conv_2_reg_33__4_ ( .D(n15206), .CK(clk), .RN(rst_n), .Q(
        conv_2[499]) );
  DFFRHQXL conv_2_reg_34__4_ ( .D(n15205), .CK(clk), .RN(rst_n), .Q(
        conv_2[514]) );
  DFFRHQXL conv_2_reg_35__4_ ( .D(n15204), .CK(clk), .RN(rst_n), .Q(
        conv_2[529]) );
  DFFRHQXL pool_reg_15__4_ ( .D(N29295), .CK(clk), .RN(rst_n), .Q(pool[79]) );
  DFFRHQXL pool_reg_17__4_ ( .D(N29305), .CK(clk), .RN(rst_n), .Q(pool[89]) );
  DFFRHQXL pool_reg_12__4_ ( .D(N29280), .CK(clk), .RN(rst_n), .Q(pool[64]) );
  DFFRHQXL pool_reg_11__4_ ( .D(N29275), .CK(clk), .RN(rst_n), .Q(pool[59]) );
  DFFRHQXL pool_reg_14__4_ ( .D(N29290), .CK(clk), .RN(rst_n), .Q(pool[74]) );
  DFFRHQXL pool_reg_9__4_ ( .D(N29265), .CK(clk), .RN(rst_n), .Q(pool[49]) );
  DFFRHQXL pool_reg_10__4_ ( .D(N29270), .CK(clk), .RN(rst_n), .Q(pool[54]) );
  DFFRHQXL pool_reg_16__4_ ( .D(N29300), .CK(clk), .RN(rst_n), .Q(pool[84]) );
  DFFRHQXL pool_reg_13__4_ ( .D(N29285), .CK(clk), .RN(rst_n), .Q(pool[69]) );
  DFFRHQXL filter_1_bias_reg_4_ ( .D(n14727), .CK(clk), .RN(rst_n), .Q(
        filter_1_bias[4]) );
  DFFRHQXL conv_1_reg_0__4_ ( .D(n16459), .CK(clk), .RN(rst_n), .Q(conv_1[4])
         );
  DFFRHQXL conv_1_reg_1__4_ ( .D(n16444), .CK(clk), .RN(rst_n), .Q(conv_1[19])
         );
  DFFRHQXL conv_1_reg_2__4_ ( .D(n16429), .CK(clk), .RN(rst_n), .Q(conv_1[34])
         );
  DFFRHQXL conv_1_reg_3__4_ ( .D(n16414), .CK(clk), .RN(rst_n), .Q(conv_1[49])
         );
  DFFRHQXL conv_1_reg_4__4_ ( .D(n16399), .CK(clk), .RN(rst_n), .Q(conv_1[64])
         );
  DFFRHQXL conv_1_reg_5__4_ ( .D(n16384), .CK(clk), .RN(rst_n), .Q(conv_1[79])
         );
  DFFRHQXL conv_1_reg_6__4_ ( .D(n16369), .CK(clk), .RN(rst_n), .Q(conv_1[94])
         );
  DFFRHQXL conv_1_reg_7__4_ ( .D(n16354), .CK(clk), .RN(rst_n), .Q(conv_1[109]) );
  DFFRHQXL conv_1_reg_8__4_ ( .D(n16339), .CK(clk), .RN(rst_n), .Q(conv_1[124]) );
  DFFRHQXL conv_1_reg_9__4_ ( .D(n16324), .CK(clk), .RN(rst_n), .Q(conv_1[139]) );
  DFFRHQXL conv_1_reg_10__4_ ( .D(n16309), .CK(clk), .RN(rst_n), .Q(
        conv_1[154]) );
  DFFRHQXL conv_1_reg_11__4_ ( .D(n16294), .CK(clk), .RN(rst_n), .Q(
        conv_1[169]) );
  DFFRHQXL conv_1_reg_12__4_ ( .D(n16279), .CK(clk), .RN(rst_n), .Q(
        conv_1[184]) );
  DFFRHQXL conv_1_reg_13__4_ ( .D(n16264), .CK(clk), .RN(rst_n), .Q(
        conv_1[199]) );
  DFFRHQXL conv_1_reg_14__4_ ( .D(n16249), .CK(clk), .RN(rst_n), .Q(
        conv_1[214]) );
  DFFRHQXL conv_1_reg_15__4_ ( .D(n16234), .CK(clk), .RN(rst_n), .Q(
        conv_1[229]) );
  DFFRHQXL conv_1_reg_16__4_ ( .D(n16219), .CK(clk), .RN(rst_n), .Q(
        conv_1[244]) );
  DFFRHQXL conv_1_reg_17__4_ ( .D(n16204), .CK(clk), .RN(rst_n), .Q(
        conv_1[259]) );
  DFFRHQXL conv_1_reg_18__4_ ( .D(n16189), .CK(clk), .RN(rst_n), .Q(
        conv_1[274]) );
  DFFRHQXL conv_1_reg_19__4_ ( .D(n16174), .CK(clk), .RN(rst_n), .Q(
        conv_1[289]) );
  DFFRHQXL conv_1_reg_20__4_ ( .D(n16159), .CK(clk), .RN(rst_n), .Q(
        conv_1[304]) );
  DFFRHQXL conv_1_reg_21__4_ ( .D(n16144), .CK(clk), .RN(rst_n), .Q(
        conv_1[319]) );
  DFFRHQXL conv_1_reg_22__4_ ( .D(n16129), .CK(clk), .RN(rst_n), .Q(
        conv_1[334]) );
  DFFRHQXL conv_1_reg_23__4_ ( .D(n16114), .CK(clk), .RN(rst_n), .Q(
        conv_1[349]) );
  DFFRHQXL conv_1_reg_24__4_ ( .D(n16099), .CK(clk), .RN(rst_n), .Q(
        conv_1[364]) );
  DFFRHQXL conv_1_reg_25__4_ ( .D(n16084), .CK(clk), .RN(rst_n), .Q(
        conv_1[379]) );
  DFFRHQXL conv_1_reg_26__4_ ( .D(n16069), .CK(clk), .RN(rst_n), .Q(
        conv_1[394]) );
  DFFRHQXL conv_1_reg_27__4_ ( .D(n16054), .CK(clk), .RN(rst_n), .Q(
        conv_1[409]) );
  DFFRHQXL conv_1_reg_28__4_ ( .D(n16039), .CK(clk), .RN(rst_n), .Q(
        conv_1[424]) );
  DFFRHQXL conv_1_reg_29__4_ ( .D(n16024), .CK(clk), .RN(rst_n), .Q(
        conv_1[439]) );
  DFFRHQXL conv_1_reg_30__4_ ( .D(n16009), .CK(clk), .RN(rst_n), .Q(
        conv_1[454]) );
  DFFRHQXL conv_1_reg_31__4_ ( .D(n15994), .CK(clk), .RN(rst_n), .Q(
        conv_1[469]) );
  DFFRHQXL conv_1_reg_32__4_ ( .D(n15979), .CK(clk), .RN(rst_n), .Q(
        conv_1[484]) );
  DFFRHQXL conv_1_reg_33__4_ ( .D(n15964), .CK(clk), .RN(rst_n), .Q(
        conv_1[499]) );
  DFFRHQXL conv_1_reg_34__4_ ( .D(n15949), .CK(clk), .RN(rst_n), .Q(
        conv_1[514]) );
  DFFRHQXL conv_1_reg_35__4_ ( .D(n15934), .CK(clk), .RN(rst_n), .Q(
        conv_1[529]) );
  DFFRHQXL pool_reg_6__4_ ( .D(N29250), .CK(clk), .RN(rst_n), .Q(pool[34]) );
  DFFRHQXL pool_reg_8__4_ ( .D(N29260), .CK(clk), .RN(rst_n), .Q(pool[44]) );
  DFFRHQXL pool_reg_3__4_ ( .D(N29235), .CK(clk), .RN(rst_n), .Q(pool[19]) );
  DFFRHQXL pool_reg_2__4_ ( .D(N29230), .CK(clk), .RN(rst_n), .Q(pool[14]) );
  DFFRHQXL pool_reg_5__4_ ( .D(N29245), .CK(clk), .RN(rst_n), .Q(pool[29]) );
  DFFRHQXL pool_reg_0__4_ ( .D(N29220), .CK(clk), .RN(rst_n), .Q(pool[4]) );
  DFFRHQXL pool_reg_1__4_ ( .D(N29225), .CK(clk), .RN(rst_n), .Q(pool[9]) );
  DFFRHQXL pool_reg_7__4_ ( .D(N29255), .CK(clk), .RN(rst_n), .Q(pool[39]) );
  DFFRHQXL pool_reg_4__4_ ( .D(N29240), .CK(clk), .RN(rst_n), .Q(pool[24]) );
  DFFRHQXL filter_3_bias_reg_3_ ( .D(n14726), .CK(clk), .RN(rst_n), .Q(
        filter_3_bias[3]) );
  DFFRHQXL conv_3_reg_0__3_ ( .D(n15815), .CK(clk), .RN(rst_n), .Q(conv_3[3])
         );
  DFFRHQXL conv_3_reg_1__3_ ( .D(n15814), .CK(clk), .RN(rst_n), .Q(conv_3[18])
         );
  DFFRHQXL conv_3_reg_2__3_ ( .D(n15813), .CK(clk), .RN(rst_n), .Q(conv_3[33])
         );
  DFFRHQXL conv_3_reg_3__3_ ( .D(n15812), .CK(clk), .RN(rst_n), .Q(conv_3[48])
         );
  DFFRHQXL conv_3_reg_4__3_ ( .D(n15811), .CK(clk), .RN(rst_n), .Q(conv_3[63])
         );
  DFFRHQXL conv_3_reg_5__3_ ( .D(n15810), .CK(clk), .RN(rst_n), .Q(conv_3[78])
         );
  DFFRHQXL conv_3_reg_6__3_ ( .D(n15809), .CK(clk), .RN(rst_n), .Q(conv_3[93])
         );
  DFFRHQXL conv_3_reg_7__3_ ( .D(n15808), .CK(clk), .RN(rst_n), .Q(conv_3[108]) );
  DFFRHQXL conv_3_reg_8__3_ ( .D(n15807), .CK(clk), .RN(rst_n), .Q(conv_3[123]) );
  DFFRHQXL conv_3_reg_9__3_ ( .D(n15806), .CK(clk), .RN(rst_n), .Q(conv_3[138]) );
  DFFRHQXL conv_3_reg_10__3_ ( .D(n15805), .CK(clk), .RN(rst_n), .Q(
        conv_3[153]) );
  DFFRHQXL conv_3_reg_11__3_ ( .D(n15804), .CK(clk), .RN(rst_n), .Q(
        conv_3[168]) );
  DFFRHQXL conv_3_reg_12__3_ ( .D(n15803), .CK(clk), .RN(rst_n), .Q(
        conv_3[183]) );
  DFFRHQXL conv_3_reg_13__3_ ( .D(n15802), .CK(clk), .RN(rst_n), .Q(
        conv_3[198]) );
  DFFRHQXL conv_3_reg_14__3_ ( .D(n15801), .CK(clk), .RN(rst_n), .Q(
        conv_3[213]) );
  DFFRHQXL conv_3_reg_15__3_ ( .D(n15800), .CK(clk), .RN(rst_n), .Q(
        conv_3[228]) );
  DFFRHQXL conv_3_reg_16__3_ ( .D(n15799), .CK(clk), .RN(rst_n), .Q(
        conv_3[243]) );
  DFFRHQXL conv_3_reg_17__3_ ( .D(n15798), .CK(clk), .RN(rst_n), .Q(
        conv_3[258]) );
  DFFRHQXL conv_3_reg_18__3_ ( .D(n15797), .CK(clk), .RN(rst_n), .Q(
        conv_3[273]) );
  DFFRHQXL conv_3_reg_19__3_ ( .D(n15796), .CK(clk), .RN(rst_n), .Q(
        conv_3[288]) );
  DFFRHQXL conv_3_reg_20__3_ ( .D(n15795), .CK(clk), .RN(rst_n), .Q(
        conv_3[303]) );
  DFFRHQXL conv_3_reg_21__3_ ( .D(n15794), .CK(clk), .RN(rst_n), .Q(
        conv_3[318]) );
  DFFRHQXL conv_3_reg_22__3_ ( .D(n15793), .CK(clk), .RN(rst_n), .Q(
        conv_3[333]) );
  DFFRHQXL conv_3_reg_23__3_ ( .D(n15792), .CK(clk), .RN(rst_n), .Q(
        conv_3[348]) );
  DFFRHQXL conv_3_reg_24__3_ ( .D(n15791), .CK(clk), .RN(rst_n), .Q(
        conv_3[363]) );
  DFFRHQXL conv_3_reg_25__3_ ( .D(n15790), .CK(clk), .RN(rst_n), .Q(
        conv_3[378]) );
  DFFRHQXL conv_3_reg_26__3_ ( .D(n15789), .CK(clk), .RN(rst_n), .Q(
        conv_3[393]) );
  DFFRHQXL conv_3_reg_27__3_ ( .D(n15788), .CK(clk), .RN(rst_n), .Q(
        conv_3[408]) );
  DFFRHQXL conv_3_reg_28__3_ ( .D(n15787), .CK(clk), .RN(rst_n), .Q(
        conv_3[423]) );
  DFFRHQXL conv_3_reg_29__3_ ( .D(n15786), .CK(clk), .RN(rst_n), .Q(
        conv_3[438]) );
  DFFRHQXL conv_3_reg_30__3_ ( .D(n15785), .CK(clk), .RN(rst_n), .Q(
        conv_3[453]) );
  DFFRHQXL conv_3_reg_31__3_ ( .D(n15784), .CK(clk), .RN(rst_n), .Q(
        conv_3[468]) );
  DFFRHQXL conv_3_reg_32__3_ ( .D(n15783), .CK(clk), .RN(rst_n), .Q(
        conv_3[483]) );
  DFFRHQXL conv_3_reg_33__3_ ( .D(n15782), .CK(clk), .RN(rst_n), .Q(
        conv_3[498]) );
  DFFRHQXL conv_3_reg_34__3_ ( .D(n15781), .CK(clk), .RN(rst_n), .Q(
        conv_3[513]) );
  DFFRHQXL conv_3_reg_35__3_ ( .D(n15780), .CK(clk), .RN(rst_n), .Q(
        conv_3[528]) );
  DFFRHQXL pool_reg_24__3_ ( .D(N29339), .CK(clk), .RN(rst_n), .Q(pool[123])
         );
  DFFRHQXL pool_reg_26__3_ ( .D(N29349), .CK(clk), .RN(rst_n), .Q(pool[133])
         );
  DFFRHQXL pool_reg_21__3_ ( .D(N29324), .CK(clk), .RN(rst_n), .Q(pool[108])
         );
  DFFRHQXL pool_reg_20__3_ ( .D(N29319), .CK(clk), .RN(rst_n), .Q(pool[103])
         );
  DFFRHQXL pool_reg_23__3_ ( .D(N29334), .CK(clk), .RN(rst_n), .Q(pool[118])
         );
  DFFRHQXL pool_reg_18__3_ ( .D(N29309), .CK(clk), .RN(rst_n), .Q(pool[93]) );
  DFFRHQXL pool_reg_19__3_ ( .D(N29314), .CK(clk), .RN(rst_n), .Q(pool[98]) );
  DFFRHQXL pool_reg_25__3_ ( .D(N29344), .CK(clk), .RN(rst_n), .Q(pool[128])
         );
  DFFRHQXL pool_reg_22__3_ ( .D(N29329), .CK(clk), .RN(rst_n), .Q(pool[113])
         );
  DFFRHQXL filter_2_bias_reg_3_ ( .D(n14725), .CK(clk), .RN(rst_n), .Q(
        filter_2_bias[3]) );
  DFFRHQXL conv_2_reg_0__3_ ( .D(n15275), .CK(clk), .RN(rst_n), .Q(conv_2[3])
         );
  DFFRHQXL conv_2_reg_1__3_ ( .D(n15274), .CK(clk), .RN(rst_n), .Q(conv_2[18])
         );
  DFFRHQXL conv_2_reg_2__3_ ( .D(n15273), .CK(clk), .RN(rst_n), .Q(conv_2[33])
         );
  DFFRHQXL conv_2_reg_3__3_ ( .D(n15272), .CK(clk), .RN(rst_n), .Q(conv_2[48])
         );
  DFFRHQXL conv_2_reg_4__3_ ( .D(n15271), .CK(clk), .RN(rst_n), .Q(conv_2[63])
         );
  DFFRHQXL conv_2_reg_5__3_ ( .D(n15270), .CK(clk), .RN(rst_n), .Q(conv_2[78])
         );
  DFFRHQXL conv_2_reg_6__3_ ( .D(n15269), .CK(clk), .RN(rst_n), .Q(conv_2[93])
         );
  DFFRHQXL conv_2_reg_7__3_ ( .D(n15268), .CK(clk), .RN(rst_n), .Q(conv_2[108]) );
  DFFRHQXL conv_2_reg_8__3_ ( .D(n15267), .CK(clk), .RN(rst_n), .Q(conv_2[123]) );
  DFFRHQXL conv_2_reg_9__3_ ( .D(n15266), .CK(clk), .RN(rst_n), .Q(conv_2[138]) );
  DFFRHQXL conv_2_reg_10__3_ ( .D(n15265), .CK(clk), .RN(rst_n), .Q(
        conv_2[153]) );
  DFFRHQXL conv_2_reg_11__3_ ( .D(n15264), .CK(clk), .RN(rst_n), .Q(
        conv_2[168]) );
  DFFRHQXL conv_2_reg_12__3_ ( .D(n15263), .CK(clk), .RN(rst_n), .Q(
        conv_2[183]) );
  DFFRHQXL conv_2_reg_13__3_ ( .D(n15262), .CK(clk), .RN(rst_n), .Q(
        conv_2[198]) );
  DFFRHQXL conv_2_reg_14__3_ ( .D(n15261), .CK(clk), .RN(rst_n), .Q(
        conv_2[213]) );
  DFFRHQXL conv_2_reg_15__3_ ( .D(n15260), .CK(clk), .RN(rst_n), .Q(
        conv_2[228]) );
  DFFRHQXL conv_2_reg_16__3_ ( .D(n15259), .CK(clk), .RN(rst_n), .Q(
        conv_2[243]) );
  DFFRHQXL conv_2_reg_17__3_ ( .D(n15258), .CK(clk), .RN(rst_n), .Q(
        conv_2[258]) );
  DFFRHQXL conv_2_reg_18__3_ ( .D(n15257), .CK(clk), .RN(rst_n), .Q(
        conv_2[273]) );
  DFFRHQXL conv_2_reg_19__3_ ( .D(n15256), .CK(clk), .RN(rst_n), .Q(
        conv_2[288]) );
  DFFRHQXL conv_2_reg_20__3_ ( .D(n15255), .CK(clk), .RN(rst_n), .Q(
        conv_2[303]) );
  DFFRHQXL conv_2_reg_21__3_ ( .D(n15254), .CK(clk), .RN(rst_n), .Q(
        conv_2[318]) );
  DFFRHQXL conv_2_reg_22__3_ ( .D(n15253), .CK(clk), .RN(rst_n), .Q(
        conv_2[333]) );
  DFFRHQXL conv_2_reg_23__3_ ( .D(n15252), .CK(clk), .RN(rst_n), .Q(
        conv_2[348]) );
  DFFRHQXL conv_2_reg_24__3_ ( .D(n15251), .CK(clk), .RN(rst_n), .Q(
        conv_2[363]) );
  DFFRHQXL conv_2_reg_25__3_ ( .D(n15250), .CK(clk), .RN(rst_n), .Q(
        conv_2[378]) );
  DFFRHQXL conv_2_reg_26__3_ ( .D(n15249), .CK(clk), .RN(rst_n), .Q(
        conv_2[393]) );
  DFFRHQXL conv_2_reg_27__3_ ( .D(n15248), .CK(clk), .RN(rst_n), .Q(
        conv_2[408]) );
  DFFRHQXL conv_2_reg_28__3_ ( .D(n15247), .CK(clk), .RN(rst_n), .Q(
        conv_2[423]) );
  DFFRHQXL conv_2_reg_29__3_ ( .D(n15246), .CK(clk), .RN(rst_n), .Q(
        conv_2[438]) );
  DFFRHQXL conv_2_reg_30__3_ ( .D(n15245), .CK(clk), .RN(rst_n), .Q(
        conv_2[453]) );
  DFFRHQXL conv_2_reg_31__3_ ( .D(n15244), .CK(clk), .RN(rst_n), .Q(
        conv_2[468]) );
  DFFRHQXL conv_2_reg_32__3_ ( .D(n15243), .CK(clk), .RN(rst_n), .Q(
        conv_2[483]) );
  DFFRHQXL conv_2_reg_33__3_ ( .D(n15242), .CK(clk), .RN(rst_n), .Q(
        conv_2[498]) );
  DFFRHQXL conv_2_reg_34__3_ ( .D(n15241), .CK(clk), .RN(rst_n), .Q(
        conv_2[513]) );
  DFFRHQXL conv_2_reg_35__3_ ( .D(n15240), .CK(clk), .RN(rst_n), .Q(
        conv_2[528]) );
  DFFRHQXL pool_reg_15__3_ ( .D(N29294), .CK(clk), .RN(rst_n), .Q(pool[78]) );
  DFFRHQXL pool_reg_17__3_ ( .D(N29304), .CK(clk), .RN(rst_n), .Q(pool[88]) );
  DFFRHQXL pool_reg_12__3_ ( .D(N29279), .CK(clk), .RN(rst_n), .Q(pool[63]) );
  DFFRHQXL pool_reg_11__3_ ( .D(N29274), .CK(clk), .RN(rst_n), .Q(pool[58]) );
  DFFRHQXL pool_reg_14__3_ ( .D(N29289), .CK(clk), .RN(rst_n), .Q(pool[73]) );
  DFFRHQXL pool_reg_9__3_ ( .D(N29264), .CK(clk), .RN(rst_n), .Q(pool[48]) );
  DFFRHQXL pool_reg_10__3_ ( .D(N29269), .CK(clk), .RN(rst_n), .Q(pool[53]) );
  DFFRHQXL pool_reg_16__3_ ( .D(N29299), .CK(clk), .RN(rst_n), .Q(pool[83]) );
  DFFRHQXL pool_reg_13__3_ ( .D(N29284), .CK(clk), .RN(rst_n), .Q(pool[68]) );
  DFFRHQXL filter_1_bias_reg_3_ ( .D(n14724), .CK(clk), .RN(rst_n), .Q(
        filter_1_bias[3]) );
  DFFRHQXL conv_1_reg_0__3_ ( .D(n16460), .CK(clk), .RN(rst_n), .Q(conv_1[3])
         );
  DFFRHQXL conv_1_reg_1__3_ ( .D(n16445), .CK(clk), .RN(rst_n), .Q(conv_1[18])
         );
  DFFRHQXL conv_1_reg_2__3_ ( .D(n16430), .CK(clk), .RN(rst_n), .Q(conv_1[33])
         );
  DFFRHQXL conv_1_reg_3__3_ ( .D(n16415), .CK(clk), .RN(rst_n), .Q(conv_1[48])
         );
  DFFRHQXL conv_1_reg_4__3_ ( .D(n16400), .CK(clk), .RN(rst_n), .Q(conv_1[63])
         );
  DFFRHQXL conv_1_reg_5__3_ ( .D(n16385), .CK(clk), .RN(rst_n), .Q(conv_1[78])
         );
  DFFRHQXL conv_1_reg_6__3_ ( .D(n16370), .CK(clk), .RN(rst_n), .Q(conv_1[93])
         );
  DFFRHQXL conv_1_reg_7__3_ ( .D(n16355), .CK(clk), .RN(rst_n), .Q(conv_1[108]) );
  DFFRHQXL conv_1_reg_8__3_ ( .D(n16340), .CK(clk), .RN(rst_n), .Q(conv_1[123]) );
  DFFRHQXL conv_1_reg_9__3_ ( .D(n16325), .CK(clk), .RN(rst_n), .Q(conv_1[138]) );
  DFFRHQXL conv_1_reg_10__3_ ( .D(n16310), .CK(clk), .RN(rst_n), .Q(
        conv_1[153]) );
  DFFRHQXL conv_1_reg_11__3_ ( .D(n16295), .CK(clk), .RN(rst_n), .Q(
        conv_1[168]) );
  DFFRHQXL conv_1_reg_12__3_ ( .D(n16280), .CK(clk), .RN(rst_n), .Q(
        conv_1[183]) );
  DFFRHQXL conv_1_reg_13__3_ ( .D(n16265), .CK(clk), .RN(rst_n), .Q(
        conv_1[198]) );
  DFFRHQXL conv_1_reg_14__3_ ( .D(n16250), .CK(clk), .RN(rst_n), .Q(
        conv_1[213]) );
  DFFRHQXL conv_1_reg_15__3_ ( .D(n16235), .CK(clk), .RN(rst_n), .Q(
        conv_1[228]) );
  DFFRHQXL conv_1_reg_16__3_ ( .D(n16220), .CK(clk), .RN(rst_n), .Q(
        conv_1[243]) );
  DFFRHQXL conv_1_reg_17__3_ ( .D(n16205), .CK(clk), .RN(rst_n), .Q(
        conv_1[258]) );
  DFFRHQXL conv_1_reg_18__3_ ( .D(n16190), .CK(clk), .RN(rst_n), .Q(
        conv_1[273]) );
  DFFRHQXL conv_1_reg_19__3_ ( .D(n16175), .CK(clk), .RN(rst_n), .Q(
        conv_1[288]) );
  DFFRHQXL conv_1_reg_20__3_ ( .D(n16160), .CK(clk), .RN(rst_n), .Q(
        conv_1[303]) );
  DFFRHQXL conv_1_reg_21__3_ ( .D(n16145), .CK(clk), .RN(rst_n), .Q(
        conv_1[318]) );
  DFFRHQXL conv_1_reg_22__3_ ( .D(n16130), .CK(clk), .RN(rst_n), .Q(
        conv_1[333]) );
  DFFRHQXL conv_1_reg_23__3_ ( .D(n16115), .CK(clk), .RN(rst_n), .Q(
        conv_1[348]) );
  DFFRHQXL conv_1_reg_24__3_ ( .D(n16100), .CK(clk), .RN(rst_n), .Q(
        conv_1[363]) );
  DFFRHQXL conv_1_reg_25__3_ ( .D(n16085), .CK(clk), .RN(rst_n), .Q(
        conv_1[378]) );
  DFFRHQXL conv_1_reg_26__3_ ( .D(n16070), .CK(clk), .RN(rst_n), .Q(
        conv_1[393]) );
  DFFRHQXL conv_1_reg_27__3_ ( .D(n16055), .CK(clk), .RN(rst_n), .Q(
        conv_1[408]) );
  DFFRHQXL conv_1_reg_28__3_ ( .D(n16040), .CK(clk), .RN(rst_n), .Q(
        conv_1[423]) );
  DFFRHQXL conv_1_reg_29__3_ ( .D(n16025), .CK(clk), .RN(rst_n), .Q(
        conv_1[438]) );
  DFFRHQXL conv_1_reg_30__3_ ( .D(n16010), .CK(clk), .RN(rst_n), .Q(
        conv_1[453]) );
  DFFRHQXL conv_1_reg_31__3_ ( .D(n15995), .CK(clk), .RN(rst_n), .Q(
        conv_1[468]) );
  DFFRHQXL conv_1_reg_32__3_ ( .D(n15980), .CK(clk), .RN(rst_n), .Q(
        conv_1[483]) );
  DFFRHQXL conv_1_reg_33__3_ ( .D(n15965), .CK(clk), .RN(rst_n), .Q(
        conv_1[498]) );
  DFFRHQXL conv_1_reg_34__3_ ( .D(n15950), .CK(clk), .RN(rst_n), .Q(
        conv_1[513]) );
  DFFRHQXL conv_1_reg_35__3_ ( .D(n15935), .CK(clk), .RN(rst_n), .Q(
        conv_1[528]) );
  DFFRHQXL pool_reg_6__3_ ( .D(N29249), .CK(clk), .RN(rst_n), .Q(pool[33]) );
  DFFRHQXL pool_reg_8__3_ ( .D(N29259), .CK(clk), .RN(rst_n), .Q(pool[43]) );
  DFFRHQXL pool_reg_3__3_ ( .D(N29234), .CK(clk), .RN(rst_n), .Q(pool[18]) );
  DFFRHQXL pool_reg_2__3_ ( .D(N29229), .CK(clk), .RN(rst_n), .Q(pool[13]) );
  DFFRHQXL pool_reg_5__3_ ( .D(N29244), .CK(clk), .RN(rst_n), .Q(pool[28]) );
  DFFRHQXL pool_reg_0__3_ ( .D(N29219), .CK(clk), .RN(rst_n), .Q(pool[3]) );
  DFFRHQXL pool_reg_1__3_ ( .D(N29224), .CK(clk), .RN(rst_n), .Q(pool[8]) );
  DFFRHQXL pool_reg_7__3_ ( .D(N29254), .CK(clk), .RN(rst_n), .Q(pool[38]) );
  DFFRHQXL pool_reg_4__3_ ( .D(N29239), .CK(clk), .RN(rst_n), .Q(pool[23]) );
  DFFRHQXL filter_3_bias_reg_2_ ( .D(n14723), .CK(clk), .RN(rst_n), .Q(
        filter_3_bias[2]) );
  DFFRHQXL conv_3_reg_0__2_ ( .D(n15851), .CK(clk), .RN(rst_n), .Q(conv_3[2])
         );
  DFFRHQXL conv_3_reg_1__2_ ( .D(n15850), .CK(clk), .RN(rst_n), .Q(conv_3[17])
         );
  DFFRHQXL conv_3_reg_2__2_ ( .D(n15849), .CK(clk), .RN(rst_n), .Q(conv_3[32])
         );
  DFFRHQXL conv_3_reg_3__2_ ( .D(n15848), .CK(clk), .RN(rst_n), .Q(conv_3[47])
         );
  DFFRHQXL conv_3_reg_4__2_ ( .D(n15847), .CK(clk), .RN(rst_n), .Q(conv_3[62])
         );
  DFFRHQXL conv_3_reg_5__2_ ( .D(n15846), .CK(clk), .RN(rst_n), .Q(conv_3[77])
         );
  DFFRHQXL conv_3_reg_6__2_ ( .D(n15845), .CK(clk), .RN(rst_n), .Q(conv_3[92])
         );
  DFFRHQXL conv_3_reg_7__2_ ( .D(n15844), .CK(clk), .RN(rst_n), .Q(conv_3[107]) );
  DFFRHQXL conv_3_reg_8__2_ ( .D(n15843), .CK(clk), .RN(rst_n), .Q(conv_3[122]) );
  DFFRHQXL conv_3_reg_9__2_ ( .D(n15842), .CK(clk), .RN(rst_n), .Q(conv_3[137]) );
  DFFRHQXL conv_3_reg_10__2_ ( .D(n15841), .CK(clk), .RN(rst_n), .Q(
        conv_3[152]) );
  DFFRHQXL conv_3_reg_11__2_ ( .D(n15840), .CK(clk), .RN(rst_n), .Q(
        conv_3[167]) );
  DFFRHQXL conv_3_reg_12__2_ ( .D(n15839), .CK(clk), .RN(rst_n), .Q(
        conv_3[182]) );
  DFFRHQXL conv_3_reg_13__2_ ( .D(n15838), .CK(clk), .RN(rst_n), .Q(
        conv_3[197]) );
  DFFRHQXL conv_3_reg_14__2_ ( .D(n15837), .CK(clk), .RN(rst_n), .Q(
        conv_3[212]) );
  DFFRHQXL conv_3_reg_15__2_ ( .D(n15836), .CK(clk), .RN(rst_n), .Q(
        conv_3[227]) );
  DFFRHQXL conv_3_reg_16__2_ ( .D(n15835), .CK(clk), .RN(rst_n), .Q(
        conv_3[242]) );
  DFFRHQXL conv_3_reg_17__2_ ( .D(n15834), .CK(clk), .RN(rst_n), .Q(
        conv_3[257]) );
  DFFRHQXL conv_3_reg_18__2_ ( .D(n15833), .CK(clk), .RN(rst_n), .Q(
        conv_3[272]) );
  DFFRHQXL conv_3_reg_19__2_ ( .D(n15832), .CK(clk), .RN(rst_n), .Q(
        conv_3[287]) );
  DFFRHQXL conv_3_reg_20__2_ ( .D(n15831), .CK(clk), .RN(rst_n), .Q(
        conv_3[302]) );
  DFFRHQXL conv_3_reg_21__2_ ( .D(n15830), .CK(clk), .RN(rst_n), .Q(
        conv_3[317]) );
  DFFRHQXL conv_3_reg_22__2_ ( .D(n15829), .CK(clk), .RN(rst_n), .Q(
        conv_3[332]) );
  DFFRHQXL conv_3_reg_23__2_ ( .D(n15828), .CK(clk), .RN(rst_n), .Q(
        conv_3[347]) );
  DFFRHQXL conv_3_reg_24__2_ ( .D(n15827), .CK(clk), .RN(rst_n), .Q(
        conv_3[362]) );
  DFFRHQXL conv_3_reg_25__2_ ( .D(n15826), .CK(clk), .RN(rst_n), .Q(
        conv_3[377]) );
  DFFRHQXL conv_3_reg_26__2_ ( .D(n15825), .CK(clk), .RN(rst_n), .Q(
        conv_3[392]) );
  DFFRHQXL conv_3_reg_27__2_ ( .D(n15824), .CK(clk), .RN(rst_n), .Q(
        conv_3[407]) );
  DFFRHQXL conv_3_reg_28__2_ ( .D(n15823), .CK(clk), .RN(rst_n), .Q(
        conv_3[422]) );
  DFFRHQXL conv_3_reg_29__2_ ( .D(n15822), .CK(clk), .RN(rst_n), .Q(
        conv_3[437]) );
  DFFRHQXL conv_3_reg_30__2_ ( .D(n15821), .CK(clk), .RN(rst_n), .Q(
        conv_3[452]) );
  DFFRHQXL conv_3_reg_31__2_ ( .D(n15820), .CK(clk), .RN(rst_n), .Q(
        conv_3[467]) );
  DFFRHQXL conv_3_reg_32__2_ ( .D(n15819), .CK(clk), .RN(rst_n), .Q(
        conv_3[482]) );
  DFFRHQXL conv_3_reg_33__2_ ( .D(n15818), .CK(clk), .RN(rst_n), .Q(
        conv_3[497]) );
  DFFRHQXL conv_3_reg_34__2_ ( .D(n15817), .CK(clk), .RN(rst_n), .Q(
        conv_3[512]) );
  DFFRHQXL conv_3_reg_35__2_ ( .D(n15816), .CK(clk), .RN(rst_n), .Q(
        conv_3[527]) );
  DFFRHQXL pool_reg_24__2_ ( .D(N29338), .CK(clk), .RN(rst_n), .Q(pool[122])
         );
  DFFRHQXL pool_reg_26__2_ ( .D(N29348), .CK(clk), .RN(rst_n), .Q(pool[132])
         );
  DFFRHQXL pool_reg_21__2_ ( .D(N29323), .CK(clk), .RN(rst_n), .Q(pool[107])
         );
  DFFRHQXL pool_reg_20__2_ ( .D(N29318), .CK(clk), .RN(rst_n), .Q(pool[102])
         );
  DFFRHQXL pool_reg_23__2_ ( .D(N29333), .CK(clk), .RN(rst_n), .Q(pool[117])
         );
  DFFRHQXL pool_reg_18__2_ ( .D(N29308), .CK(clk), .RN(rst_n), .Q(pool[92]) );
  DFFRHQXL pool_reg_19__2_ ( .D(N29313), .CK(clk), .RN(rst_n), .Q(pool[97]) );
  DFFRHQXL pool_reg_25__2_ ( .D(N29343), .CK(clk), .RN(rst_n), .Q(pool[127])
         );
  DFFRHQXL pool_reg_22__2_ ( .D(N29328), .CK(clk), .RN(rst_n), .Q(pool[112])
         );
  DFFRHQXL filter_2_bias_reg_2_ ( .D(n14722), .CK(clk), .RN(rst_n), .Q(
        filter_2_bias[2]) );
  DFFRHQXL conv_2_reg_0__2_ ( .D(n15311), .CK(clk), .RN(rst_n), .Q(conv_2[2])
         );
  DFFRHQXL conv_2_reg_1__2_ ( .D(n15310), .CK(clk), .RN(rst_n), .Q(conv_2[17])
         );
  DFFRHQXL conv_2_reg_2__2_ ( .D(n15309), .CK(clk), .RN(rst_n), .Q(conv_2[32])
         );
  DFFRHQXL conv_2_reg_3__2_ ( .D(n15308), .CK(clk), .RN(rst_n), .Q(conv_2[47])
         );
  DFFRHQXL conv_2_reg_4__2_ ( .D(n15307), .CK(clk), .RN(rst_n), .Q(conv_2[62])
         );
  DFFRHQXL conv_2_reg_5__2_ ( .D(n15306), .CK(clk), .RN(rst_n), .Q(conv_2[77])
         );
  DFFRHQXL conv_2_reg_6__2_ ( .D(n15305), .CK(clk), .RN(rst_n), .Q(conv_2[92])
         );
  DFFRHQXL conv_2_reg_7__2_ ( .D(n15304), .CK(clk), .RN(rst_n), .Q(conv_2[107]) );
  DFFRHQXL conv_2_reg_8__2_ ( .D(n15303), .CK(clk), .RN(rst_n), .Q(conv_2[122]) );
  DFFRHQXL conv_2_reg_9__2_ ( .D(n15302), .CK(clk), .RN(rst_n), .Q(conv_2[137]) );
  DFFRHQXL conv_2_reg_10__2_ ( .D(n15301), .CK(clk), .RN(rst_n), .Q(
        conv_2[152]) );
  DFFRHQXL conv_2_reg_11__2_ ( .D(n15300), .CK(clk), .RN(rst_n), .Q(
        conv_2[167]) );
  DFFRHQXL conv_2_reg_12__2_ ( .D(n15299), .CK(clk), .RN(rst_n), .Q(
        conv_2[182]) );
  DFFRHQXL conv_2_reg_13__2_ ( .D(n15298), .CK(clk), .RN(rst_n), .Q(
        conv_2[197]) );
  DFFRHQXL conv_2_reg_14__2_ ( .D(n15297), .CK(clk), .RN(rst_n), .Q(
        conv_2[212]) );
  DFFRHQXL conv_2_reg_15__2_ ( .D(n15296), .CK(clk), .RN(rst_n), .Q(
        conv_2[227]) );
  DFFRHQXL conv_2_reg_16__2_ ( .D(n15295), .CK(clk), .RN(rst_n), .Q(
        conv_2[242]) );
  DFFRHQXL conv_2_reg_17__2_ ( .D(n15294), .CK(clk), .RN(rst_n), .Q(
        conv_2[257]) );
  DFFRHQXL conv_2_reg_18__2_ ( .D(n15293), .CK(clk), .RN(rst_n), .Q(
        conv_2[272]) );
  DFFRHQXL conv_2_reg_19__2_ ( .D(n15292), .CK(clk), .RN(rst_n), .Q(
        conv_2[287]) );
  DFFRHQXL conv_2_reg_20__2_ ( .D(n15291), .CK(clk), .RN(rst_n), .Q(
        conv_2[302]) );
  DFFRHQXL conv_2_reg_21__2_ ( .D(n15290), .CK(clk), .RN(rst_n), .Q(
        conv_2[317]) );
  DFFRHQXL conv_2_reg_22__2_ ( .D(n15289), .CK(clk), .RN(rst_n), .Q(
        conv_2[332]) );
  DFFRHQXL conv_2_reg_23__2_ ( .D(n15288), .CK(clk), .RN(rst_n), .Q(
        conv_2[347]) );
  DFFRHQXL conv_2_reg_24__2_ ( .D(n15287), .CK(clk), .RN(rst_n), .Q(
        conv_2[362]) );
  DFFRHQXL conv_2_reg_25__2_ ( .D(n15286), .CK(clk), .RN(rst_n), .Q(
        conv_2[377]) );
  DFFRHQXL conv_2_reg_26__2_ ( .D(n15285), .CK(clk), .RN(rst_n), .Q(
        conv_2[392]) );
  DFFRHQXL conv_2_reg_27__2_ ( .D(n15284), .CK(clk), .RN(rst_n), .Q(
        conv_2[407]) );
  DFFRHQXL conv_2_reg_28__2_ ( .D(n15283), .CK(clk), .RN(rst_n), .Q(
        conv_2[422]) );
  DFFRHQXL conv_2_reg_29__2_ ( .D(n15282), .CK(clk), .RN(rst_n), .Q(
        conv_2[437]) );
  DFFRHQXL conv_2_reg_30__2_ ( .D(n15281), .CK(clk), .RN(rst_n), .Q(
        conv_2[452]) );
  DFFRHQXL conv_2_reg_31__2_ ( .D(n15280), .CK(clk), .RN(rst_n), .Q(
        conv_2[467]) );
  DFFRHQXL conv_2_reg_32__2_ ( .D(n15279), .CK(clk), .RN(rst_n), .Q(
        conv_2[482]) );
  DFFRHQXL conv_2_reg_33__2_ ( .D(n15278), .CK(clk), .RN(rst_n), .Q(
        conv_2[497]) );
  DFFRHQXL conv_2_reg_34__2_ ( .D(n15277), .CK(clk), .RN(rst_n), .Q(
        conv_2[512]) );
  DFFRHQXL conv_2_reg_35__2_ ( .D(n15276), .CK(clk), .RN(rst_n), .Q(
        conv_2[527]) );
  DFFRHQXL pool_reg_15__2_ ( .D(N29293), .CK(clk), .RN(rst_n), .Q(pool[77]) );
  DFFRHQXL pool_reg_17__2_ ( .D(N29303), .CK(clk), .RN(rst_n), .Q(pool[87]) );
  DFFRHQXL pool_reg_12__2_ ( .D(N29278), .CK(clk), .RN(rst_n), .Q(pool[62]) );
  DFFRHQXL pool_reg_11__2_ ( .D(N29273), .CK(clk), .RN(rst_n), .Q(pool[57]) );
  DFFRHQXL pool_reg_14__2_ ( .D(N29288), .CK(clk), .RN(rst_n), .Q(pool[72]) );
  DFFRHQXL pool_reg_9__2_ ( .D(N29263), .CK(clk), .RN(rst_n), .Q(pool[47]) );
  DFFRHQXL pool_reg_10__2_ ( .D(N29268), .CK(clk), .RN(rst_n), .Q(pool[52]) );
  DFFRHQXL pool_reg_16__2_ ( .D(N29298), .CK(clk), .RN(rst_n), .Q(pool[82]) );
  DFFRHQXL pool_reg_13__2_ ( .D(N29283), .CK(clk), .RN(rst_n), .Q(pool[67]) );
  DFFRHQXL filter_1_bias_reg_2_ ( .D(n14721), .CK(clk), .RN(rst_n), .Q(
        filter_1_bias[2]) );
  DFFRHQXL conv_1_reg_0__2_ ( .D(n16461), .CK(clk), .RN(rst_n), .Q(conv_1[2])
         );
  DFFRHQXL conv_1_reg_1__2_ ( .D(n16446), .CK(clk), .RN(rst_n), .Q(conv_1[17])
         );
  DFFRHQXL conv_1_reg_2__2_ ( .D(n16431), .CK(clk), .RN(rst_n), .Q(conv_1[32])
         );
  DFFRHQXL conv_1_reg_3__2_ ( .D(n16416), .CK(clk), .RN(rst_n), .Q(conv_1[47])
         );
  DFFRHQXL conv_1_reg_4__2_ ( .D(n16401), .CK(clk), .RN(rst_n), .Q(conv_1[62])
         );
  DFFRHQXL conv_1_reg_5__2_ ( .D(n16386), .CK(clk), .RN(rst_n), .Q(conv_1[77])
         );
  DFFRHQXL conv_1_reg_6__2_ ( .D(n16371), .CK(clk), .RN(rst_n), .Q(conv_1[92])
         );
  DFFRHQXL conv_1_reg_7__2_ ( .D(n16356), .CK(clk), .RN(rst_n), .Q(conv_1[107]) );
  DFFRHQXL conv_1_reg_8__2_ ( .D(n16341), .CK(clk), .RN(rst_n), .Q(conv_1[122]) );
  DFFRHQXL conv_1_reg_9__2_ ( .D(n16326), .CK(clk), .RN(rst_n), .Q(conv_1[137]) );
  DFFRHQXL conv_1_reg_10__2_ ( .D(n16311), .CK(clk), .RN(rst_n), .Q(
        conv_1[152]) );
  DFFRHQXL conv_1_reg_11__2_ ( .D(n16296), .CK(clk), .RN(rst_n), .Q(
        conv_1[167]) );
  DFFRHQXL conv_1_reg_12__2_ ( .D(n16281), .CK(clk), .RN(rst_n), .Q(
        conv_1[182]) );
  DFFRHQXL conv_1_reg_13__2_ ( .D(n16266), .CK(clk), .RN(rst_n), .Q(
        conv_1[197]) );
  DFFRHQXL conv_1_reg_14__2_ ( .D(n16251), .CK(clk), .RN(rst_n), .Q(
        conv_1[212]) );
  DFFRHQXL conv_1_reg_15__2_ ( .D(n16236), .CK(clk), .RN(rst_n), .Q(
        conv_1[227]) );
  DFFRHQXL conv_1_reg_16__2_ ( .D(n16221), .CK(clk), .RN(rst_n), .Q(
        conv_1[242]) );
  DFFRHQXL conv_1_reg_17__2_ ( .D(n16206), .CK(clk), .RN(rst_n), .Q(
        conv_1[257]) );
  DFFRHQXL conv_1_reg_18__2_ ( .D(n16191), .CK(clk), .RN(rst_n), .Q(
        conv_1[272]) );
  DFFRHQXL conv_1_reg_19__2_ ( .D(n16176), .CK(clk), .RN(rst_n), .Q(
        conv_1[287]) );
  DFFRHQXL conv_1_reg_20__2_ ( .D(n16161), .CK(clk), .RN(rst_n), .Q(
        conv_1[302]) );
  DFFRHQXL conv_1_reg_21__2_ ( .D(n16146), .CK(clk), .RN(rst_n), .Q(
        conv_1[317]) );
  DFFRHQXL conv_1_reg_22__2_ ( .D(n16131), .CK(clk), .RN(rst_n), .Q(
        conv_1[332]) );
  DFFRHQXL conv_1_reg_23__2_ ( .D(n16116), .CK(clk), .RN(rst_n), .Q(
        conv_1[347]) );
  DFFRHQXL conv_1_reg_24__2_ ( .D(n16101), .CK(clk), .RN(rst_n), .Q(
        conv_1[362]) );
  DFFRHQXL conv_1_reg_25__2_ ( .D(n16086), .CK(clk), .RN(rst_n), .Q(
        conv_1[377]) );
  DFFRHQXL conv_1_reg_26__2_ ( .D(n16071), .CK(clk), .RN(rst_n), .Q(
        conv_1[392]) );
  DFFRHQXL conv_1_reg_27__2_ ( .D(n16056), .CK(clk), .RN(rst_n), .Q(
        conv_1[407]) );
  DFFRHQXL conv_1_reg_28__2_ ( .D(n16041), .CK(clk), .RN(rst_n), .Q(
        conv_1[422]) );
  DFFRHQXL conv_1_reg_29__2_ ( .D(n16026), .CK(clk), .RN(rst_n), .Q(
        conv_1[437]) );
  DFFRHQXL conv_1_reg_30__2_ ( .D(n16011), .CK(clk), .RN(rst_n), .Q(
        conv_1[452]) );
  DFFRHQXL conv_1_reg_31__2_ ( .D(n15996), .CK(clk), .RN(rst_n), .Q(
        conv_1[467]) );
  DFFRHQXL conv_1_reg_32__2_ ( .D(n15981), .CK(clk), .RN(rst_n), .Q(
        conv_1[482]) );
  DFFRHQXL conv_1_reg_33__2_ ( .D(n15966), .CK(clk), .RN(rst_n), .Q(
        conv_1[497]) );
  DFFRHQXL conv_1_reg_34__2_ ( .D(n15951), .CK(clk), .RN(rst_n), .Q(
        conv_1[512]) );
  DFFRHQXL conv_1_reg_35__2_ ( .D(n15936), .CK(clk), .RN(rst_n), .Q(
        conv_1[527]) );
  DFFRHQXL pool_reg_6__2_ ( .D(N29248), .CK(clk), .RN(rst_n), .Q(pool[32]) );
  DFFRHQXL pool_reg_8__2_ ( .D(N29258), .CK(clk), .RN(rst_n), .Q(pool[42]) );
  DFFRHQXL pool_reg_3__2_ ( .D(N29233), .CK(clk), .RN(rst_n), .Q(pool[17]) );
  DFFRHQXL pool_reg_2__2_ ( .D(N29228), .CK(clk), .RN(rst_n), .Q(pool[12]) );
  DFFRHQXL pool_reg_5__2_ ( .D(N29243), .CK(clk), .RN(rst_n), .Q(pool[27]) );
  DFFRHQXL pool_reg_0__2_ ( .D(N29218), .CK(clk), .RN(rst_n), .Q(pool[2]) );
  DFFRHQXL pool_reg_1__2_ ( .D(N29223), .CK(clk), .RN(rst_n), .Q(pool[7]) );
  DFFRHQXL pool_reg_7__2_ ( .D(N29253), .CK(clk), .RN(rst_n), .Q(pool[37]) );
  DFFRHQXL pool_reg_4__2_ ( .D(N29238), .CK(clk), .RN(rst_n), .Q(pool[22]) );
  DFFRHQXL filter_3_bias_reg_1_ ( .D(n14720), .CK(clk), .RN(rst_n), .Q(
        filter_3_bias[1]) );
  DFFRHQXL conv_3_reg_0__1_ ( .D(n15887), .CK(clk), .RN(rst_n), .Q(conv_3[1])
         );
  DFFRHQXL conv_3_reg_1__1_ ( .D(n15886), .CK(clk), .RN(rst_n), .Q(conv_3[16])
         );
  DFFRHQXL conv_3_reg_2__1_ ( .D(n15885), .CK(clk), .RN(rst_n), .Q(conv_3[31])
         );
  DFFRHQXL conv_3_reg_3__1_ ( .D(n15884), .CK(clk), .RN(rst_n), .Q(conv_3[46])
         );
  DFFRHQXL conv_3_reg_4__1_ ( .D(n15883), .CK(clk), .RN(rst_n), .Q(conv_3[61])
         );
  DFFRHQXL conv_3_reg_5__1_ ( .D(n15882), .CK(clk), .RN(rst_n), .Q(conv_3[76])
         );
  DFFRHQXL conv_3_reg_6__1_ ( .D(n15881), .CK(clk), .RN(rst_n), .Q(conv_3[91])
         );
  DFFRHQXL conv_3_reg_7__1_ ( .D(n15880), .CK(clk), .RN(rst_n), .Q(conv_3[106]) );
  DFFRHQXL conv_3_reg_8__1_ ( .D(n15879), .CK(clk), .RN(rst_n), .Q(conv_3[121]) );
  DFFRHQXL conv_3_reg_9__1_ ( .D(n15878), .CK(clk), .RN(rst_n), .Q(conv_3[136]) );
  DFFRHQXL conv_3_reg_10__1_ ( .D(n15877), .CK(clk), .RN(rst_n), .Q(
        conv_3[151]) );
  DFFRHQXL conv_3_reg_11__1_ ( .D(n15876), .CK(clk), .RN(rst_n), .Q(
        conv_3[166]) );
  DFFRHQXL conv_3_reg_12__1_ ( .D(n15875), .CK(clk), .RN(rst_n), .Q(
        conv_3[181]) );
  DFFRHQXL conv_3_reg_13__1_ ( .D(n15874), .CK(clk), .RN(rst_n), .Q(
        conv_3[196]) );
  DFFRHQXL conv_3_reg_14__1_ ( .D(n15873), .CK(clk), .RN(rst_n), .Q(
        conv_3[211]) );
  DFFRHQXL conv_3_reg_15__1_ ( .D(n15872), .CK(clk), .RN(rst_n), .Q(
        conv_3[226]) );
  DFFRHQXL conv_3_reg_16__1_ ( .D(n15871), .CK(clk), .RN(rst_n), .Q(
        conv_3[241]) );
  DFFRHQXL conv_3_reg_17__1_ ( .D(n15870), .CK(clk), .RN(rst_n), .Q(
        conv_3[256]) );
  DFFRHQXL conv_3_reg_18__1_ ( .D(n15869), .CK(clk), .RN(rst_n), .Q(
        conv_3[271]) );
  DFFRHQXL conv_3_reg_19__1_ ( .D(n15868), .CK(clk), .RN(rst_n), .Q(
        conv_3[286]) );
  DFFRHQXL conv_3_reg_20__1_ ( .D(n15867), .CK(clk), .RN(rst_n), .Q(
        conv_3[301]) );
  DFFRHQXL conv_3_reg_21__1_ ( .D(n15866), .CK(clk), .RN(rst_n), .Q(
        conv_3[316]) );
  DFFRHQXL conv_3_reg_22__1_ ( .D(n15865), .CK(clk), .RN(rst_n), .Q(
        conv_3[331]) );
  DFFRHQXL conv_3_reg_23__1_ ( .D(n15864), .CK(clk), .RN(rst_n), .Q(
        conv_3[346]) );
  DFFRHQXL conv_3_reg_24__1_ ( .D(n15863), .CK(clk), .RN(rst_n), .Q(
        conv_3[361]) );
  DFFRHQXL conv_3_reg_25__1_ ( .D(n15862), .CK(clk), .RN(rst_n), .Q(
        conv_3[376]) );
  DFFRHQXL conv_3_reg_26__1_ ( .D(n15861), .CK(clk), .RN(rst_n), .Q(
        conv_3[391]) );
  DFFRHQXL conv_3_reg_27__1_ ( .D(n15860), .CK(clk), .RN(rst_n), .Q(
        conv_3[406]) );
  DFFRHQXL conv_3_reg_28__1_ ( .D(n15859), .CK(clk), .RN(rst_n), .Q(
        conv_3[421]) );
  DFFRHQXL conv_3_reg_29__1_ ( .D(n15858), .CK(clk), .RN(rst_n), .Q(
        conv_3[436]) );
  DFFRHQXL conv_3_reg_30__1_ ( .D(n15857), .CK(clk), .RN(rst_n), .Q(
        conv_3[451]) );
  DFFRHQXL conv_3_reg_31__1_ ( .D(n15856), .CK(clk), .RN(rst_n), .Q(
        conv_3[466]) );
  DFFRHQXL conv_3_reg_32__1_ ( .D(n15855), .CK(clk), .RN(rst_n), .Q(
        conv_3[481]) );
  DFFRHQXL conv_3_reg_33__1_ ( .D(n15854), .CK(clk), .RN(rst_n), .Q(
        conv_3[496]) );
  DFFRHQXL conv_3_reg_34__1_ ( .D(n15853), .CK(clk), .RN(rst_n), .Q(
        conv_3[511]) );
  DFFRHQXL conv_3_reg_35__1_ ( .D(n15852), .CK(clk), .RN(rst_n), .Q(
        conv_3[526]) );
  DFFRHQXL pool_reg_24__1_ ( .D(N29337), .CK(clk), .RN(rst_n), .Q(pool[121])
         );
  DFFRHQXL pool_reg_26__1_ ( .D(N29347), .CK(clk), .RN(rst_n), .Q(pool[131])
         );
  DFFRHQXL pool_reg_21__1_ ( .D(N29322), .CK(clk), .RN(rst_n), .Q(pool[106])
         );
  DFFRHQXL pool_reg_20__1_ ( .D(N29317), .CK(clk), .RN(rst_n), .Q(pool[101])
         );
  DFFRHQXL pool_reg_23__1_ ( .D(N29332), .CK(clk), .RN(rst_n), .Q(pool[116])
         );
  DFFRHQXL pool_reg_18__1_ ( .D(N29307), .CK(clk), .RN(rst_n), .Q(pool[91]) );
  DFFRHQXL pool_reg_19__1_ ( .D(N29312), .CK(clk), .RN(rst_n), .Q(pool[96]) );
  DFFRHQXL pool_reg_25__1_ ( .D(N29342), .CK(clk), .RN(rst_n), .Q(pool[126])
         );
  DFFRHQXL pool_reg_22__1_ ( .D(N29327), .CK(clk), .RN(rst_n), .Q(pool[111])
         );
  DFFRHQXL filter_2_bias_reg_1_ ( .D(n14719), .CK(clk), .RN(rst_n), .Q(
        filter_2_bias[1]) );
  DFFRHQXL conv_2_reg_0__1_ ( .D(n15347), .CK(clk), .RN(rst_n), .Q(conv_2[1])
         );
  DFFRHQXL conv_2_reg_1__1_ ( .D(n15346), .CK(clk), .RN(rst_n), .Q(conv_2[16])
         );
  DFFRHQXL conv_2_reg_2__1_ ( .D(n15345), .CK(clk), .RN(rst_n), .Q(conv_2[31])
         );
  DFFRHQXL conv_2_reg_3__1_ ( .D(n15344), .CK(clk), .RN(rst_n), .Q(conv_2[46])
         );
  DFFRHQXL conv_2_reg_4__1_ ( .D(n15343), .CK(clk), .RN(rst_n), .Q(conv_2[61])
         );
  DFFRHQXL conv_2_reg_5__1_ ( .D(n15342), .CK(clk), .RN(rst_n), .Q(conv_2[76])
         );
  DFFRHQXL conv_2_reg_6__1_ ( .D(n15341), .CK(clk), .RN(rst_n), .Q(conv_2[91])
         );
  DFFRHQXL conv_2_reg_7__1_ ( .D(n15340), .CK(clk), .RN(rst_n), .Q(conv_2[106]) );
  DFFRHQXL conv_2_reg_8__1_ ( .D(n15339), .CK(clk), .RN(rst_n), .Q(conv_2[121]) );
  DFFRHQXL conv_2_reg_9__1_ ( .D(n15338), .CK(clk), .RN(rst_n), .Q(conv_2[136]) );
  DFFRHQXL conv_2_reg_10__1_ ( .D(n15337), .CK(clk), .RN(rst_n), .Q(
        conv_2[151]) );
  DFFRHQXL conv_2_reg_11__1_ ( .D(n15336), .CK(clk), .RN(rst_n), .Q(
        conv_2[166]) );
  DFFRHQXL conv_2_reg_12__1_ ( .D(n15335), .CK(clk), .RN(rst_n), .Q(
        conv_2[181]) );
  DFFRHQXL conv_2_reg_13__1_ ( .D(n15334), .CK(clk), .RN(rst_n), .Q(
        conv_2[196]) );
  DFFRHQXL conv_2_reg_14__1_ ( .D(n15333), .CK(clk), .RN(rst_n), .Q(
        conv_2[211]) );
  DFFRHQXL conv_2_reg_15__1_ ( .D(n15332), .CK(clk), .RN(rst_n), .Q(
        conv_2[226]) );
  DFFRHQXL conv_2_reg_16__1_ ( .D(n15331), .CK(clk), .RN(rst_n), .Q(
        conv_2[241]) );
  DFFRHQXL conv_2_reg_17__1_ ( .D(n15330), .CK(clk), .RN(rst_n), .Q(
        conv_2[256]) );
  DFFRHQXL conv_2_reg_18__1_ ( .D(n15329), .CK(clk), .RN(rst_n), .Q(
        conv_2[271]) );
  DFFRHQXL conv_2_reg_19__1_ ( .D(n15328), .CK(clk), .RN(rst_n), .Q(
        conv_2[286]) );
  DFFRHQXL conv_2_reg_20__1_ ( .D(n15327), .CK(clk), .RN(rst_n), .Q(
        conv_2[301]) );
  DFFRHQXL conv_2_reg_21__1_ ( .D(n15326), .CK(clk), .RN(rst_n), .Q(
        conv_2[316]) );
  DFFRHQXL conv_2_reg_22__1_ ( .D(n15325), .CK(clk), .RN(rst_n), .Q(
        conv_2[331]) );
  DFFRHQXL conv_2_reg_23__1_ ( .D(n15324), .CK(clk), .RN(rst_n), .Q(
        conv_2[346]) );
  DFFRHQXL conv_2_reg_24__1_ ( .D(n15323), .CK(clk), .RN(rst_n), .Q(
        conv_2[361]) );
  DFFRHQXL conv_2_reg_25__1_ ( .D(n15322), .CK(clk), .RN(rst_n), .Q(
        conv_2[376]) );
  DFFRHQXL conv_2_reg_26__1_ ( .D(n15321), .CK(clk), .RN(rst_n), .Q(
        conv_2[391]) );
  DFFRHQXL conv_2_reg_27__1_ ( .D(n15320), .CK(clk), .RN(rst_n), .Q(
        conv_2[406]) );
  DFFRHQXL conv_2_reg_28__1_ ( .D(n15319), .CK(clk), .RN(rst_n), .Q(
        conv_2[421]) );
  DFFRHQXL conv_2_reg_29__1_ ( .D(n15318), .CK(clk), .RN(rst_n), .Q(
        conv_2[436]) );
  DFFRHQXL conv_2_reg_30__1_ ( .D(n15317), .CK(clk), .RN(rst_n), .Q(
        conv_2[451]) );
  DFFRHQXL conv_2_reg_31__1_ ( .D(n15316), .CK(clk), .RN(rst_n), .Q(
        conv_2[466]) );
  DFFRHQXL conv_2_reg_32__1_ ( .D(n15315), .CK(clk), .RN(rst_n), .Q(
        conv_2[481]) );
  DFFRHQXL conv_2_reg_33__1_ ( .D(n15314), .CK(clk), .RN(rst_n), .Q(
        conv_2[496]) );
  DFFRHQXL conv_2_reg_34__1_ ( .D(n15313), .CK(clk), .RN(rst_n), .Q(
        conv_2[511]) );
  DFFRHQXL conv_2_reg_35__1_ ( .D(n15312), .CK(clk), .RN(rst_n), .Q(
        conv_2[526]) );
  DFFRHQXL pool_reg_15__1_ ( .D(N29292), .CK(clk), .RN(rst_n), .Q(pool[76]) );
  DFFRHQXL pool_reg_17__1_ ( .D(N29302), .CK(clk), .RN(rst_n), .Q(pool[86]) );
  DFFRHQXL pool_reg_12__1_ ( .D(N29277), .CK(clk), .RN(rst_n), .Q(pool[61]) );
  DFFRHQXL pool_reg_11__1_ ( .D(N29272), .CK(clk), .RN(rst_n), .Q(pool[56]) );
  DFFRHQXL pool_reg_14__1_ ( .D(N29287), .CK(clk), .RN(rst_n), .Q(pool[71]) );
  DFFRHQXL pool_reg_9__1_ ( .D(N29262), .CK(clk), .RN(rst_n), .Q(pool[46]) );
  DFFRHQXL pool_reg_10__1_ ( .D(N29267), .CK(clk), .RN(rst_n), .Q(pool[51]) );
  DFFRHQXL pool_reg_16__1_ ( .D(N29297), .CK(clk), .RN(rst_n), .Q(pool[81]) );
  DFFRHQXL pool_reg_13__1_ ( .D(N29282), .CK(clk), .RN(rst_n), .Q(pool[66]) );
  DFFRHQXL filter_1_bias_reg_1_ ( .D(n14718), .CK(clk), .RN(rst_n), .Q(
        filter_1_bias[1]) );
  DFFRHQXL conv_1_reg_0__1_ ( .D(n16462), .CK(clk), .RN(rst_n), .Q(conv_1[1])
         );
  DFFRHQXL conv_1_reg_1__1_ ( .D(n16447), .CK(clk), .RN(rst_n), .Q(conv_1[16])
         );
  DFFRHQXL conv_1_reg_2__1_ ( .D(n16432), .CK(clk), .RN(rst_n), .Q(conv_1[31])
         );
  DFFRHQXL conv_1_reg_3__1_ ( .D(n16417), .CK(clk), .RN(rst_n), .Q(conv_1[46])
         );
  DFFRHQXL conv_1_reg_4__1_ ( .D(n16402), .CK(clk), .RN(rst_n), .Q(conv_1[61])
         );
  DFFRHQXL conv_1_reg_5__1_ ( .D(n16387), .CK(clk), .RN(rst_n), .Q(conv_1[76])
         );
  DFFRHQXL conv_1_reg_6__1_ ( .D(n16372), .CK(clk), .RN(rst_n), .Q(conv_1[91])
         );
  DFFRHQXL conv_1_reg_7__1_ ( .D(n16357), .CK(clk), .RN(rst_n), .Q(conv_1[106]) );
  DFFRHQXL conv_1_reg_8__1_ ( .D(n16342), .CK(clk), .RN(rst_n), .Q(conv_1[121]) );
  DFFRHQXL conv_1_reg_9__1_ ( .D(n16327), .CK(clk), .RN(rst_n), .Q(conv_1[136]) );
  DFFRHQXL conv_1_reg_10__1_ ( .D(n16312), .CK(clk), .RN(rst_n), .Q(
        conv_1[151]) );
  DFFRHQXL conv_1_reg_11__1_ ( .D(n16297), .CK(clk), .RN(rst_n), .Q(
        conv_1[166]) );
  DFFRHQXL conv_1_reg_12__1_ ( .D(n16282), .CK(clk), .RN(rst_n), .Q(
        conv_1[181]) );
  DFFRHQXL conv_1_reg_13__1_ ( .D(n16267), .CK(clk), .RN(rst_n), .Q(
        conv_1[196]) );
  DFFRHQXL conv_1_reg_14__1_ ( .D(n16252), .CK(clk), .RN(rst_n), .Q(
        conv_1[211]) );
  DFFRHQXL conv_1_reg_15__1_ ( .D(n16237), .CK(clk), .RN(rst_n), .Q(
        conv_1[226]) );
  DFFRHQXL conv_1_reg_16__1_ ( .D(n16222), .CK(clk), .RN(rst_n), .Q(
        conv_1[241]) );
  DFFRHQXL conv_1_reg_17__1_ ( .D(n16207), .CK(clk), .RN(rst_n), .Q(
        conv_1[256]) );
  DFFRHQXL conv_1_reg_18__1_ ( .D(n16192), .CK(clk), .RN(rst_n), .Q(
        conv_1[271]) );
  DFFRHQXL conv_1_reg_19__1_ ( .D(n16177), .CK(clk), .RN(rst_n), .Q(
        conv_1[286]) );
  DFFRHQXL conv_1_reg_20__1_ ( .D(n16162), .CK(clk), .RN(rst_n), .Q(
        conv_1[301]) );
  DFFRHQXL conv_1_reg_21__1_ ( .D(n16147), .CK(clk), .RN(rst_n), .Q(
        conv_1[316]) );
  DFFRHQXL conv_1_reg_22__1_ ( .D(n16132), .CK(clk), .RN(rst_n), .Q(
        conv_1[331]) );
  DFFRHQXL conv_1_reg_23__1_ ( .D(n16117), .CK(clk), .RN(rst_n), .Q(
        conv_1[346]) );
  DFFRHQXL conv_1_reg_24__1_ ( .D(n16102), .CK(clk), .RN(rst_n), .Q(
        conv_1[361]) );
  DFFRHQXL conv_1_reg_25__1_ ( .D(n16087), .CK(clk), .RN(rst_n), .Q(
        conv_1[376]) );
  DFFRHQXL conv_1_reg_26__1_ ( .D(n16072), .CK(clk), .RN(rst_n), .Q(
        conv_1[391]) );
  DFFRHQXL conv_1_reg_27__1_ ( .D(n16057), .CK(clk), .RN(rst_n), .Q(
        conv_1[406]) );
  DFFRHQXL conv_1_reg_28__1_ ( .D(n16042), .CK(clk), .RN(rst_n), .Q(
        conv_1[421]) );
  DFFRHQXL conv_1_reg_29__1_ ( .D(n16027), .CK(clk), .RN(rst_n), .Q(
        conv_1[436]) );
  DFFRHQXL conv_1_reg_30__1_ ( .D(n16012), .CK(clk), .RN(rst_n), .Q(
        conv_1[451]) );
  DFFRHQXL conv_1_reg_31__1_ ( .D(n15997), .CK(clk), .RN(rst_n), .Q(
        conv_1[466]) );
  DFFRHQXL conv_1_reg_32__1_ ( .D(n15982), .CK(clk), .RN(rst_n), .Q(
        conv_1[481]) );
  DFFRHQXL conv_1_reg_33__1_ ( .D(n15967), .CK(clk), .RN(rst_n), .Q(
        conv_1[496]) );
  DFFRHQXL conv_1_reg_34__1_ ( .D(n15952), .CK(clk), .RN(rst_n), .Q(
        conv_1[511]) );
  DFFRHQXL conv_1_reg_35__1_ ( .D(n15937), .CK(clk), .RN(rst_n), .Q(
        conv_1[526]) );
  DFFRHQXL pool_reg_6__1_ ( .D(N29247), .CK(clk), .RN(rst_n), .Q(pool[31]) );
  DFFRHQXL pool_reg_8__1_ ( .D(N29257), .CK(clk), .RN(rst_n), .Q(pool[41]) );
  DFFRHQXL pool_reg_3__1_ ( .D(N29232), .CK(clk), .RN(rst_n), .Q(pool[16]) );
  DFFRHQXL pool_reg_2__1_ ( .D(N29227), .CK(clk), .RN(rst_n), .Q(pool[11]) );
  DFFRHQXL pool_reg_5__1_ ( .D(N29242), .CK(clk), .RN(rst_n), .Q(pool[26]) );
  DFFRHQXL pool_reg_0__1_ ( .D(N29217), .CK(clk), .RN(rst_n), .Q(pool[1]) );
  DFFRHQXL pool_reg_1__1_ ( .D(N29222), .CK(clk), .RN(rst_n), .Q(pool[6]) );
  DFFRHQXL pool_reg_7__1_ ( .D(N29252), .CK(clk), .RN(rst_n), .Q(pool[36]) );
  DFFRHQXL pool_reg_4__1_ ( .D(N29237), .CK(clk), .RN(rst_n), .Q(pool[21]) );
  DFFRHQXL filter_1_reg_8__0_ ( .D(n14717), .CK(clk), .RN(rst_n), .Q(
        filter_1[48]) );
  DFFRHQXL filter_1_reg_7__0_ ( .D(n14716), .CK(clk), .RN(rst_n), .Q(
        filter_1[42]) );
  DFFRHQXL filter_1_reg_6__0_ ( .D(n14715), .CK(clk), .RN(rst_n), .Q(
        filter_1[36]) );
  DFFRHQXL filter_1_reg_5__0_ ( .D(n14714), .CK(clk), .RN(rst_n), .Q(
        filter_1[30]) );
  DFFRHQXL filter_1_reg_4__0_ ( .D(n14713), .CK(clk), .RN(rst_n), .Q(
        filter_1[24]) );
  DFFRHQXL filter_1_reg_3__0_ ( .D(n14712), .CK(clk), .RN(rst_n), .Q(
        filter_1[18]) );
  DFFRHQXL filter_1_reg_2__0_ ( .D(n14711), .CK(clk), .RN(rst_n), .Q(
        filter_1[12]) );
  DFFRHQXL filter_1_reg_1__0_ ( .D(n14710), .CK(clk), .RN(rst_n), .Q(
        filter_1[6]) );
  DFFRHQXL filter_1_reg_0__0_ ( .D(n14709), .CK(clk), .RN(rst_n), .Q(
        filter_1[0]) );
  DFFRHQXL filter_1_reg_8__1_ ( .D(n14708), .CK(clk), .RN(rst_n), .Q(
        filter_1[49]) );
  DFFRHQXL filter_1_reg_7__1_ ( .D(n14707), .CK(clk), .RN(rst_n), .Q(
        filter_1[43]) );
  DFFRHQXL filter_1_reg_6__1_ ( .D(n14706), .CK(clk), .RN(rst_n), .Q(
        filter_1[37]) );
  DFFRHQXL filter_1_reg_5__1_ ( .D(n14705), .CK(clk), .RN(rst_n), .Q(
        filter_1[31]) );
  DFFRHQXL filter_1_reg_4__1_ ( .D(n14704), .CK(clk), .RN(rst_n), .Q(
        filter_1[25]) );
  DFFRHQXL filter_1_reg_3__1_ ( .D(n14703), .CK(clk), .RN(rst_n), .Q(
        filter_1[19]) );
  DFFRHQXL filter_1_reg_2__1_ ( .D(n14702), .CK(clk), .RN(rst_n), .Q(
        filter_1[13]) );
  DFFRHQXL filter_1_reg_1__1_ ( .D(n14701), .CK(clk), .RN(rst_n), .Q(
        filter_1[7]) );
  DFFRHQXL filter_1_reg_0__1_ ( .D(n14700), .CK(clk), .RN(rst_n), .Q(
        filter_1[1]) );
  DFFRHQXL filter_1_reg_8__2_ ( .D(n14699), .CK(clk), .RN(rst_n), .Q(
        filter_1[50]) );
  DFFRHQXL filter_1_reg_7__2_ ( .D(n14698), .CK(clk), .RN(rst_n), .Q(
        filter_1[44]) );
  DFFRHQXL filter_1_reg_6__2_ ( .D(n14697), .CK(clk), .RN(rst_n), .Q(
        filter_1[38]) );
  DFFRHQXL filter_1_reg_5__2_ ( .D(n14696), .CK(clk), .RN(rst_n), .Q(
        filter_1[32]) );
  DFFRHQXL filter_1_reg_4__2_ ( .D(n14695), .CK(clk), .RN(rst_n), .Q(
        filter_1[26]) );
  DFFRHQXL filter_1_reg_3__2_ ( .D(n14694), .CK(clk), .RN(rst_n), .Q(
        filter_1[20]) );
  DFFRHQXL filter_1_reg_2__2_ ( .D(n14693), .CK(clk), .RN(rst_n), .Q(
        filter_1[14]) );
  DFFRHQXL filter_1_reg_1__2_ ( .D(n14692), .CK(clk), .RN(rst_n), .Q(
        filter_1[8]) );
  DFFRHQXL filter_1_reg_0__2_ ( .D(n14691), .CK(clk), .RN(rst_n), .Q(
        filter_1[2]) );
  DFFRHQXL filter_1_reg_8__3_ ( .D(n14690), .CK(clk), .RN(rst_n), .Q(
        filter_1[51]) );
  DFFRHQXL filter_1_reg_7__3_ ( .D(n14689), .CK(clk), .RN(rst_n), .Q(
        filter_1[45]) );
  DFFRHQXL filter_1_reg_6__3_ ( .D(n14688), .CK(clk), .RN(rst_n), .Q(
        filter_1[39]) );
  DFFRHQXL filter_1_reg_5__3_ ( .D(n14687), .CK(clk), .RN(rst_n), .Q(
        filter_1[33]) );
  DFFRHQXL filter_1_reg_4__3_ ( .D(n14686), .CK(clk), .RN(rst_n), .Q(
        filter_1[27]) );
  DFFRHQXL filter_1_reg_3__3_ ( .D(n14685), .CK(clk), .RN(rst_n), .Q(
        filter_1[21]) );
  DFFRHQXL filter_1_reg_2__3_ ( .D(n14684), .CK(clk), .RN(rst_n), .Q(
        filter_1[15]) );
  DFFRHQXL filter_1_reg_1__3_ ( .D(n14683), .CK(clk), .RN(rst_n), .Q(
        filter_1[9]) );
  DFFRHQXL filter_1_reg_0__3_ ( .D(n14682), .CK(clk), .RN(rst_n), .Q(
        filter_1[3]) );
  DFFRHQXL filter_1_reg_8__4_ ( .D(n14681), .CK(clk), .RN(rst_n), .Q(
        filter_1[52]) );
  DFFRHQXL filter_1_reg_7__4_ ( .D(n14680), .CK(clk), .RN(rst_n), .Q(
        filter_1[46]) );
  DFFRHQXL filter_1_reg_6__4_ ( .D(n14679), .CK(clk), .RN(rst_n), .Q(
        filter_1[40]) );
  DFFRHQXL filter_1_reg_5__4_ ( .D(n14678), .CK(clk), .RN(rst_n), .Q(
        filter_1[34]) );
  DFFRHQXL filter_1_reg_4__4_ ( .D(n14677), .CK(clk), .RN(rst_n), .Q(
        filter_1[28]) );
  DFFRHQXL filter_1_reg_3__4_ ( .D(n14676), .CK(clk), .RN(rst_n), .Q(
        filter_1[22]) );
  DFFRHQXL filter_1_reg_2__4_ ( .D(n14675), .CK(clk), .RN(rst_n), .Q(
        filter_1[16]) );
  DFFRHQXL filter_1_reg_1__4_ ( .D(n14674), .CK(clk), .RN(rst_n), .Q(
        filter_1[10]) );
  DFFRHQXL filter_1_reg_0__4_ ( .D(n14673), .CK(clk), .RN(rst_n), .Q(
        filter_1[4]) );
  DFFRHQXL filter_1_reg_8__5_ ( .D(n14672), .CK(clk), .RN(rst_n), .Q(
        filter_1[53]) );
  DFFRHQXL filter_1_reg_7__5_ ( .D(n14671), .CK(clk), .RN(rst_n), .Q(
        filter_1[47]) );
  DFFRHQXL filter_1_reg_6__5_ ( .D(n14670), .CK(clk), .RN(rst_n), .Q(
        filter_1[41]) );
  DFFRHQXL filter_1_reg_5__5_ ( .D(n14669), .CK(clk), .RN(rst_n), .Q(
        filter_1[35]) );
  DFFRHQXL filter_1_reg_4__5_ ( .D(n14668), .CK(clk), .RN(rst_n), .Q(
        filter_1[29]) );
  DFFRHQXL filter_1_reg_3__5_ ( .D(n14667), .CK(clk), .RN(rst_n), .Q(
        filter_1[23]) );
  DFFRHQXL filter_1_reg_2__5_ ( .D(n14666), .CK(clk), .RN(rst_n), .Q(
        filter_1[17]) );
  DFFRHQXL filter_1_reg_1__5_ ( .D(n14665), .CK(clk), .RN(rst_n), .Q(
        filter_1[11]) );
  DFFRHQXL filter_1_reg_0__5_ ( .D(n14664), .CK(clk), .RN(rst_n), .Q(
        filter_1[5]) );
  DFFRHQXL weight_2_bias_3_reg_0_ ( .D(n14663), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_3[0]) );
  DFFRHQXL affine_2_reg_2__0_ ( .D(n16561), .CK(clk), .RN(rst_n), .Q(
        affine_2[32]) );
  DFFRHQXL weight_2_bias_2_reg_0_ ( .D(n14662), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_2[0]) );
  DFFRHQXL affine_2_reg_1__0_ ( .D(n16545), .CK(clk), .RN(rst_n), .Q(
        affine_2[16]) );
  DFFRHQXL weight_2_bias_1_reg_0_ ( .D(n14661), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_1[0]) );
  DFFRHQXL affine_2_reg_0__0_ ( .D(n16579), .CK(clk), .RN(rst_n), .Q(
        affine_2[0]) );
  DFFRHQXL weight_2_bias_3_reg_5_ ( .D(n14660), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_3[5]) );
  DFFRHQXL affine_2_reg_2__5_ ( .D(n16556), .CK(clk), .RN(rst_n), .Q(
        affine_2[37]) );
  DFFRHQXL affine_2_reg_2__6_ ( .D(n16555), .CK(clk), .RN(rst_n), .Q(
        affine_2[38]) );
  DFFRHQXL affine_2_reg_2__7_ ( .D(n16554), .CK(clk), .RN(rst_n), .Q(
        affine_2[39]) );
  DFFRHQXL affine_2_reg_2__8_ ( .D(n16553), .CK(clk), .RN(rst_n), .Q(
        affine_2[40]) );
  DFFRHQXL affine_2_reg_2__9_ ( .D(n16552), .CK(clk), .RN(rst_n), .Q(
        affine_2[41]) );
  DFFRHQXL affine_2_reg_2__10_ ( .D(n16551), .CK(clk), .RN(rst_n), .Q(
        affine_2[42]) );
  DFFRHQXL affine_2_reg_2__11_ ( .D(n16550), .CK(clk), .RN(rst_n), .Q(
        affine_2[43]) );
  DFFRHQXL affine_2_reg_2__12_ ( .D(n16549), .CK(clk), .RN(rst_n), .Q(
        affine_2[44]) );
  DFFRHQXL affine_2_reg_2__13_ ( .D(n16548), .CK(clk), .RN(rst_n), .Q(
        affine_2[45]) );
  DFFRHQXL affine_2_reg_2__14_ ( .D(n16547), .CK(clk), .RN(rst_n), .Q(
        affine_2[46]) );
  DFFRHQXL affine_2_reg_2__15_ ( .D(n16546), .CK(clk), .RN(rst_n), .Q(
        affine_2[47]) );
  DFFRHQXL weight_2_bias_2_reg_5_ ( .D(n14659), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_2[5]) );
  DFFRHQXL affine_2_reg_1__5_ ( .D(n16540), .CK(clk), .RN(rst_n), .Q(
        affine_2[21]) );
  DFFRHQXL affine_2_reg_1__6_ ( .D(n16539), .CK(clk), .RN(rst_n), .Q(
        affine_2[22]) );
  DFFRHQXL affine_2_reg_1__7_ ( .D(n16538), .CK(clk), .RN(rst_n), .Q(
        affine_2[23]) );
  DFFRHQXL affine_2_reg_1__8_ ( .D(n16537), .CK(clk), .RN(rst_n), .Q(
        affine_2[24]) );
  DFFRHQXL affine_2_reg_1__9_ ( .D(n16536), .CK(clk), .RN(rst_n), .Q(
        affine_2[25]) );
  DFFRHQXL affine_2_reg_1__10_ ( .D(n16535), .CK(clk), .RN(rst_n), .Q(
        affine_2[26]) );
  DFFRHQXL affine_2_reg_1__11_ ( .D(n16534), .CK(clk), .RN(rst_n), .Q(
        affine_2[27]) );
  DFFRHQXL affine_2_reg_1__12_ ( .D(n16533), .CK(clk), .RN(rst_n), .Q(
        affine_2[28]) );
  DFFRHQXL affine_2_reg_1__13_ ( .D(n16532), .CK(clk), .RN(rst_n), .Q(
        affine_2[29]) );
  DFFRHQXL affine_2_reg_1__14_ ( .D(n16531), .CK(clk), .RN(rst_n), .Q(
        affine_2[30]) );
  DFFRHQXL affine_2_reg_1__15_ ( .D(n16530), .CK(clk), .RN(rst_n), .Q(
        affine_2[31]) );
  DFFRHQXL weight_2_bias_1_reg_5_ ( .D(n14658), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_1[5]) );
  DFFRHQXL affine_2_reg_0__5_ ( .D(n16574), .CK(clk), .RN(rst_n), .Q(
        affine_2[5]) );
  DFFRHQXL affine_2_reg_0__6_ ( .D(n16573), .CK(clk), .RN(rst_n), .Q(
        affine_2[6]) );
  DFFRHQXL affine_2_reg_0__7_ ( .D(n16572), .CK(clk), .RN(rst_n), .Q(
        affine_2[7]) );
  DFFRHQXL affine_2_reg_0__8_ ( .D(n16571), .CK(clk), .RN(rst_n), .Q(
        affine_2[8]) );
  DFFRHQXL affine_2_reg_0__9_ ( .D(n16570), .CK(clk), .RN(rst_n), .Q(
        affine_2[9]) );
  DFFRHQXL affine_2_reg_0__10_ ( .D(n16569), .CK(clk), .RN(rst_n), .Q(
        affine_2[10]) );
  DFFRHQXL affine_2_reg_0__11_ ( .D(n16568), .CK(clk), .RN(rst_n), .Q(
        affine_2[11]) );
  DFFRHQXL affine_2_reg_0__12_ ( .D(n16567), .CK(clk), .RN(rst_n), .Q(
        affine_2[12]) );
  DFFRHQXL affine_2_reg_0__13_ ( .D(n16566), .CK(clk), .RN(rst_n), .Q(
        affine_2[13]) );
  DFFRHQXL affine_2_reg_0__14_ ( .D(n16565), .CK(clk), .RN(rst_n), .Q(
        affine_2[14]) );
  DFFRHQXL affine_2_reg_0__15_ ( .D(n16564), .CK(clk), .RN(rst_n), .Q(
        affine_2[15]) );
  DFFRHQXL weight_2_bias_3_reg_4_ ( .D(n14657), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_3[4]) );
  DFFRHQXL affine_2_reg_2__4_ ( .D(n16557), .CK(clk), .RN(rst_n), .Q(
        affine_2[36]) );
  DFFRHQXL weight_2_bias_2_reg_4_ ( .D(n14656), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_2[4]) );
  DFFRHQXL affine_2_reg_1__4_ ( .D(n16541), .CK(clk), .RN(rst_n), .Q(
        affine_2[20]) );
  DFFRHQXL weight_2_bias_1_reg_4_ ( .D(n14655), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_1[4]) );
  DFFRHQXL affine_2_reg_0__4_ ( .D(n16575), .CK(clk), .RN(rst_n), .Q(
        affine_2[4]) );
  DFFRHQXL weight_2_bias_3_reg_3_ ( .D(n14654), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_3[3]) );
  DFFRHQXL affine_2_reg_2__3_ ( .D(n16558), .CK(clk), .RN(rst_n), .Q(
        affine_2[35]) );
  DFFRHQXL weight_2_bias_2_reg_3_ ( .D(n14653), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_2[3]) );
  DFFRHQXL affine_2_reg_1__3_ ( .D(n16542), .CK(clk), .RN(rst_n), .Q(
        affine_2[19]) );
  DFFRHQXL weight_2_bias_1_reg_3_ ( .D(n14652), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_1[3]) );
  DFFRHQXL affine_2_reg_0__3_ ( .D(n16576), .CK(clk), .RN(rst_n), .Q(
        affine_2[3]) );
  DFFRHQXL weight_2_bias_3_reg_2_ ( .D(n14651), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_3[2]) );
  DFFRHQXL affine_2_reg_2__2_ ( .D(n16559), .CK(clk), .RN(rst_n), .Q(
        affine_2[34]) );
  DFFRHQXL weight_2_bias_2_reg_2_ ( .D(n14650), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_2[2]) );
  DFFRHQXL affine_2_reg_1__2_ ( .D(n16543), .CK(clk), .RN(rst_n), .Q(
        affine_2[18]) );
  DFFRHQXL weight_2_bias_1_reg_2_ ( .D(n14649), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_1[2]) );
  DFFRHQXL affine_2_reg_0__2_ ( .D(n16577), .CK(clk), .RN(rst_n), .Q(
        affine_2[2]) );
  DFFRHQXL weight_2_bias_3_reg_1_ ( .D(n14648), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_3[1]) );
  DFFRHQXL affine_2_reg_2__1_ ( .D(n16560), .CK(clk), .RN(rst_n), .Q(
        affine_2[33]) );
  DFFRHQXL weight_2_bias_2_reg_1_ ( .D(n14647), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_2[1]) );
  DFFRHQXL affine_2_reg_1__1_ ( .D(n16544), .CK(clk), .RN(rst_n), .Q(
        affine_2[17]) );
  DFFRHQXL weight_2_bias_1_reg_1_ ( .D(n14646), .CK(clk), .RN(rst_n), .Q(
        weight_2_bias_1[1]) );
  DFFRHQXL affine_2_reg_0__1_ ( .D(n16578), .CK(clk), .RN(rst_n), .Q(
        affine_2[1]) );
  DFFRHQXL weight_2_reg_8__0_ ( .D(n14645), .CK(clk), .RN(rst_n), .Q(
        weight_2[48]) );
  DFFRHQXL weight_2_reg_7__0_ ( .D(n14644), .CK(clk), .RN(rst_n), .Q(
        weight_2[42]) );
  DFFRHQXL weight_2_reg_6__0_ ( .D(n14643), .CK(clk), .RN(rst_n), .Q(
        weight_2[36]) );
  DFFRHQXL weight_2_reg_5__0_ ( .D(n14642), .CK(clk), .RN(rst_n), .Q(
        weight_2[30]) );
  DFFRHQXL weight_2_reg_4__0_ ( .D(n14641), .CK(clk), .RN(rst_n), .Q(
        weight_2[24]) );
  DFFRHQXL weight_2_reg_3__0_ ( .D(n14640), .CK(clk), .RN(rst_n), .Q(
        weight_2[18]) );
  DFFRHQXL weight_2_reg_2__0_ ( .D(n14639), .CK(clk), .RN(rst_n), .Q(
        weight_2[12]) );
  DFFRHQXL weight_2_reg_1__0_ ( .D(n14638), .CK(clk), .RN(rst_n), .Q(
        weight_2[6]) );
  DFFRHQXL weight_2_reg_0__0_ ( .D(n14637), .CK(clk), .RN(rst_n), .Q(
        weight_2[0]) );
  DFFRHQXL weight_2_reg_8__1_ ( .D(n14636), .CK(clk), .RN(rst_n), .Q(
        weight_2[49]) );
  DFFRHQXL weight_2_reg_7__1_ ( .D(n14635), .CK(clk), .RN(rst_n), .Q(
        weight_2[43]) );
  DFFRHQXL weight_2_reg_6__1_ ( .D(n14634), .CK(clk), .RN(rst_n), .Q(
        weight_2[37]) );
  DFFRHQXL weight_2_reg_5__1_ ( .D(n14633), .CK(clk), .RN(rst_n), .Q(
        weight_2[31]) );
  DFFRHQXL weight_2_reg_4__1_ ( .D(n14632), .CK(clk), .RN(rst_n), .Q(
        weight_2[25]) );
  DFFRHQXL weight_2_reg_3__1_ ( .D(n14631), .CK(clk), .RN(rst_n), .Q(
        weight_2[19]) );
  DFFRHQXL weight_2_reg_2__1_ ( .D(n14630), .CK(clk), .RN(rst_n), .Q(
        weight_2[13]) );
  DFFRHQXL weight_2_reg_1__1_ ( .D(n14629), .CK(clk), .RN(rst_n), .Q(
        weight_2[7]) );
  DFFRHQXL weight_2_reg_0__1_ ( .D(n14628), .CK(clk), .RN(rst_n), .Q(
        weight_2[1]) );
  DFFRHQXL weight_2_reg_8__2_ ( .D(n14627), .CK(clk), .RN(rst_n), .Q(
        weight_2[50]) );
  DFFRHQXL weight_2_reg_7__2_ ( .D(n14626), .CK(clk), .RN(rst_n), .Q(
        weight_2[44]) );
  DFFRHQXL weight_2_reg_6__2_ ( .D(n14625), .CK(clk), .RN(rst_n), .Q(
        weight_2[38]) );
  DFFRHQXL weight_2_reg_5__2_ ( .D(n14624), .CK(clk), .RN(rst_n), .Q(
        weight_2[32]) );
  DFFRHQXL weight_2_reg_4__2_ ( .D(n14623), .CK(clk), .RN(rst_n), .Q(
        weight_2[26]) );
  DFFRHQXL weight_2_reg_3__2_ ( .D(n14622), .CK(clk), .RN(rst_n), .Q(
        weight_2[20]) );
  DFFRHQXL weight_2_reg_2__2_ ( .D(n14621), .CK(clk), .RN(rst_n), .Q(
        weight_2[14]) );
  DFFRHQXL weight_2_reg_1__2_ ( .D(n14620), .CK(clk), .RN(rst_n), .Q(
        weight_2[8]) );
  DFFRHQXL weight_2_reg_0__2_ ( .D(n14619), .CK(clk), .RN(rst_n), .Q(
        weight_2[2]) );
  DFFRHQXL weight_2_reg_8__3_ ( .D(n14618), .CK(clk), .RN(rst_n), .Q(
        weight_2[51]) );
  DFFRHQXL weight_2_reg_7__3_ ( .D(n14617), .CK(clk), .RN(rst_n), .Q(
        weight_2[45]) );
  DFFRHQXL weight_2_reg_6__3_ ( .D(n14616), .CK(clk), .RN(rst_n), .Q(
        weight_2[39]) );
  DFFRHQXL weight_2_reg_5__3_ ( .D(n14615), .CK(clk), .RN(rst_n), .Q(
        weight_2[33]) );
  DFFRHQXL weight_2_reg_4__3_ ( .D(n14614), .CK(clk), .RN(rst_n), .Q(
        weight_2[27]) );
  DFFRHQXL weight_2_reg_3__3_ ( .D(n14613), .CK(clk), .RN(rst_n), .Q(
        weight_2[21]) );
  DFFRHQXL weight_2_reg_2__3_ ( .D(n14612), .CK(clk), .RN(rst_n), .Q(
        weight_2[15]) );
  DFFRHQXL weight_2_reg_1__3_ ( .D(n14611), .CK(clk), .RN(rst_n), .Q(
        weight_2[9]) );
  DFFRHQXL weight_2_reg_0__3_ ( .D(n14610), .CK(clk), .RN(rst_n), .Q(
        weight_2[3]) );
  DFFRHQXL weight_2_reg_8__4_ ( .D(n14609), .CK(clk), .RN(rst_n), .Q(
        weight_2[52]) );
  DFFRHQXL weight_2_reg_7__4_ ( .D(n14608), .CK(clk), .RN(rst_n), .Q(
        weight_2[46]) );
  DFFRHQXL weight_2_reg_6__4_ ( .D(n14607), .CK(clk), .RN(rst_n), .Q(
        weight_2[40]) );
  DFFRHQXL weight_2_reg_5__4_ ( .D(n14606), .CK(clk), .RN(rst_n), .Q(
        weight_2[34]) );
  DFFRHQXL weight_2_reg_4__4_ ( .D(n14605), .CK(clk), .RN(rst_n), .Q(
        weight_2[28]) );
  DFFRHQXL weight_2_reg_3__4_ ( .D(n14604), .CK(clk), .RN(rst_n), .Q(
        weight_2[22]) );
  DFFRHQXL weight_2_reg_2__4_ ( .D(n14603), .CK(clk), .RN(rst_n), .Q(
        weight_2[16]) );
  DFFRHQXL weight_2_reg_1__4_ ( .D(n14602), .CK(clk), .RN(rst_n), .Q(
        weight_2[10]) );
  DFFRHQXL weight_2_reg_0__4_ ( .D(n14601), .CK(clk), .RN(rst_n), .Q(
        weight_2[4]) );
  DFFRHQXL weight_2_reg_8__5_ ( .D(n14600), .CK(clk), .RN(rst_n), .Q(
        weight_2[53]) );
  DFFRHQXL weight_2_reg_7__5_ ( .D(n14599), .CK(clk), .RN(rst_n), .Q(
        weight_2[47]) );
  DFFRHQXL weight_2_reg_6__5_ ( .D(n14598), .CK(clk), .RN(rst_n), .Q(
        weight_2[41]) );
  DFFRHQXL weight_2_reg_5__5_ ( .D(n14597), .CK(clk), .RN(rst_n), .Q(
        weight_2[35]) );
  DFFRHQXL weight_2_reg_4__5_ ( .D(n14596), .CK(clk), .RN(rst_n), .Q(
        weight_2[29]) );
  DFFRHQXL weight_2_reg_3__5_ ( .D(n14595), .CK(clk), .RN(rst_n), .Q(
        weight_2[23]) );
  DFFRHQXL weight_2_reg_2__5_ ( .D(n14594), .CK(clk), .RN(rst_n), .Q(
        weight_2[17]) );
  DFFRHQXL weight_2_reg_1__5_ ( .D(n14593), .CK(clk), .RN(rst_n), .Q(
        weight_2[11]) );
  DFFRHQXL weight_2_reg_0__5_ ( .D(n14592), .CK(clk), .RN(rst_n), .Q(
        weight_2[5]) );
  DFFRHQXL weight_1_reg_80__0_ ( .D(n14591), .CK(clk), .RN(rst_n), .Q(
        weight_1[480]) );
  DFFRHQXL weight_1_reg_79__0_ ( .D(n14590), .CK(clk), .RN(rst_n), .Q(
        weight_1[474]) );
  DFFRHQXL weight_1_reg_78__0_ ( .D(n14589), .CK(clk), .RN(rst_n), .Q(
        weight_1[468]) );
  DFFRHQXL weight_1_reg_77__0_ ( .D(n14588), .CK(clk), .RN(rst_n), .Q(
        weight_1[462]) );
  DFFRHQXL weight_1_reg_76__0_ ( .D(n14587), .CK(clk), .RN(rst_n), .Q(
        weight_1[456]) );
  DFFRHQXL weight_1_reg_75__0_ ( .D(n14586), .CK(clk), .RN(rst_n), .Q(
        weight_1[450]) );
  DFFRHQXL weight_1_reg_74__0_ ( .D(n14585), .CK(clk), .RN(rst_n), .Q(
        weight_1[444]) );
  DFFRHQXL weight_1_reg_73__0_ ( .D(n14584), .CK(clk), .RN(rst_n), .Q(
        weight_1[438]) );
  DFFRHQXL weight_1_reg_72__0_ ( .D(n14583), .CK(clk), .RN(rst_n), .Q(
        weight_1[432]) );
  DFFRHQXL weight_1_reg_71__0_ ( .D(n14582), .CK(clk), .RN(rst_n), .Q(
        weight_1[426]) );
  DFFRHQXL weight_1_reg_70__0_ ( .D(n14581), .CK(clk), .RN(rst_n), .Q(
        weight_1[420]) );
  DFFRHQXL weight_1_reg_69__0_ ( .D(n14580), .CK(clk), .RN(rst_n), .Q(
        weight_1[414]) );
  DFFRHQXL weight_1_reg_68__0_ ( .D(n14579), .CK(clk), .RN(rst_n), .Q(
        weight_1[408]) );
  DFFRHQXL weight_1_reg_67__0_ ( .D(n14578), .CK(clk), .RN(rst_n), .Q(
        weight_1[402]) );
  DFFRHQXL weight_1_reg_66__0_ ( .D(n14577), .CK(clk), .RN(rst_n), .Q(
        weight_1[396]) );
  DFFRHQXL weight_1_reg_65__0_ ( .D(n14576), .CK(clk), .RN(rst_n), .Q(
        weight_1[390]) );
  DFFRHQXL weight_1_reg_64__0_ ( .D(n14575), .CK(clk), .RN(rst_n), .Q(
        weight_1[384]) );
  DFFRHQXL weight_1_reg_63__0_ ( .D(n14574), .CK(clk), .RN(rst_n), .Q(
        weight_1[378]) );
  DFFRHQXL weight_1_reg_62__0_ ( .D(n14573), .CK(clk), .RN(rst_n), .Q(
        weight_1[372]) );
  DFFRHQXL weight_1_reg_61__0_ ( .D(n14572), .CK(clk), .RN(rst_n), .Q(
        weight_1[366]) );
  DFFRHQXL weight_1_reg_60__0_ ( .D(n14571), .CK(clk), .RN(rst_n), .Q(
        weight_1[360]) );
  DFFRHQXL weight_1_reg_59__0_ ( .D(n14570), .CK(clk), .RN(rst_n), .Q(
        weight_1[354]) );
  DFFRHQXL weight_1_reg_58__0_ ( .D(n14569), .CK(clk), .RN(rst_n), .Q(
        weight_1[348]) );
  DFFRHQXL weight_1_reg_57__0_ ( .D(n14568), .CK(clk), .RN(rst_n), .Q(
        weight_1[342]) );
  DFFRHQXL weight_1_reg_56__0_ ( .D(n14567), .CK(clk), .RN(rst_n), .Q(
        weight_1[336]) );
  DFFRHQXL weight_1_reg_55__0_ ( .D(n14566), .CK(clk), .RN(rst_n), .Q(
        weight_1[330]) );
  DFFRHQXL weight_1_reg_54__0_ ( .D(n14565), .CK(clk), .RN(rst_n), .Q(
        weight_1[324]) );
  DFFRHQXL weight_1_reg_53__0_ ( .D(n14564), .CK(clk), .RN(rst_n), .Q(
        weight_1[318]) );
  DFFRHQXL weight_1_reg_52__0_ ( .D(n14563), .CK(clk), .RN(rst_n), .Q(
        weight_1[312]) );
  DFFRHQXL weight_1_reg_51__0_ ( .D(n14562), .CK(clk), .RN(rst_n), .Q(
        weight_1[306]) );
  DFFRHQXL weight_1_reg_50__0_ ( .D(n14561), .CK(clk), .RN(rst_n), .Q(
        weight_1[300]) );
  DFFRHQXL weight_1_reg_49__0_ ( .D(n14560), .CK(clk), .RN(rst_n), .Q(
        weight_1[294]) );
  DFFRHQXL weight_1_reg_48__0_ ( .D(n14559), .CK(clk), .RN(rst_n), .Q(
        weight_1[288]) );
  DFFRHQXL weight_1_reg_47__0_ ( .D(n14558), .CK(clk), .RN(rst_n), .Q(
        weight_1[282]) );
  DFFRHQXL weight_1_reg_46__0_ ( .D(n14557), .CK(clk), .RN(rst_n), .Q(
        weight_1[276]) );
  DFFRHQXL weight_1_reg_45__0_ ( .D(n14556), .CK(clk), .RN(rst_n), .Q(
        weight_1[270]) );
  DFFRHQXL weight_1_reg_44__0_ ( .D(n14555), .CK(clk), .RN(rst_n), .Q(
        weight_1[264]) );
  DFFRHQXL weight_1_reg_43__0_ ( .D(n14554), .CK(clk), .RN(rst_n), .Q(
        weight_1[258]) );
  DFFRHQXL weight_1_reg_42__0_ ( .D(n14553), .CK(clk), .RN(rst_n), .Q(
        weight_1[252]) );
  DFFRHQXL weight_1_reg_41__0_ ( .D(n14552), .CK(clk), .RN(rst_n), .Q(
        weight_1[246]) );
  DFFRHQXL weight_1_reg_40__0_ ( .D(n14551), .CK(clk), .RN(rst_n), .Q(
        weight_1[240]) );
  DFFRHQXL weight_1_reg_39__0_ ( .D(n14550), .CK(clk), .RN(rst_n), .Q(
        weight_1[234]) );
  DFFRHQXL weight_1_reg_38__0_ ( .D(n14549), .CK(clk), .RN(rst_n), .Q(
        weight_1[228]) );
  DFFRHQXL weight_1_reg_37__0_ ( .D(n14548), .CK(clk), .RN(rst_n), .Q(
        weight_1[222]) );
  DFFRHQXL weight_1_reg_36__0_ ( .D(n14547), .CK(clk), .RN(rst_n), .Q(
        weight_1[216]) );
  DFFRHQXL weight_1_reg_35__0_ ( .D(n14546), .CK(clk), .RN(rst_n), .Q(
        weight_1[210]) );
  DFFRHQXL weight_1_reg_34__0_ ( .D(n14545), .CK(clk), .RN(rst_n), .Q(
        weight_1[204]) );
  DFFRHQXL weight_1_reg_33__0_ ( .D(n14544), .CK(clk), .RN(rst_n), .Q(
        weight_1[198]) );
  DFFRHQXL weight_1_reg_32__0_ ( .D(n14543), .CK(clk), .RN(rst_n), .Q(
        weight_1[192]) );
  DFFRHQXL weight_1_reg_31__0_ ( .D(n14542), .CK(clk), .RN(rst_n), .Q(
        weight_1[186]) );
  DFFRHQXL weight_1_reg_30__0_ ( .D(n14541), .CK(clk), .RN(rst_n), .Q(
        weight_1[180]) );
  DFFRHQXL weight_1_reg_29__0_ ( .D(n14540), .CK(clk), .RN(rst_n), .Q(
        weight_1[174]) );
  DFFRHQXL weight_1_reg_28__0_ ( .D(n14539), .CK(clk), .RN(rst_n), .Q(
        weight_1[168]) );
  DFFRHQXL weight_1_reg_27__0_ ( .D(n14538), .CK(clk), .RN(rst_n), .Q(
        weight_1[162]) );
  DFFRHQXL weight_1_reg_26__0_ ( .D(n14537), .CK(clk), .RN(rst_n), .Q(
        weight_1[156]) );
  DFFRHQXL weight_1_reg_25__0_ ( .D(n14536), .CK(clk), .RN(rst_n), .Q(
        weight_1[150]) );
  DFFRHQXL weight_1_reg_24__0_ ( .D(n14535), .CK(clk), .RN(rst_n), .Q(
        weight_1[144]) );
  DFFRHQXL weight_1_reg_23__0_ ( .D(n14534), .CK(clk), .RN(rst_n), .Q(
        weight_1[138]) );
  DFFRHQXL weight_1_reg_22__0_ ( .D(n14533), .CK(clk), .RN(rst_n), .Q(
        weight_1[132]) );
  DFFRHQXL weight_1_reg_21__0_ ( .D(n14532), .CK(clk), .RN(rst_n), .Q(
        weight_1[126]) );
  DFFRHQXL weight_1_reg_20__0_ ( .D(n14531), .CK(clk), .RN(rst_n), .Q(
        weight_1[120]) );
  DFFRHQXL weight_1_reg_19__0_ ( .D(n14530), .CK(clk), .RN(rst_n), .Q(
        weight_1[114]) );
  DFFRHQXL weight_1_reg_18__0_ ( .D(n14529), .CK(clk), .RN(rst_n), .Q(
        weight_1[108]) );
  DFFRHQXL weight_1_reg_17__0_ ( .D(n14528), .CK(clk), .RN(rst_n), .Q(
        weight_1[102]) );
  DFFRHQXL weight_1_reg_16__0_ ( .D(n14527), .CK(clk), .RN(rst_n), .Q(
        weight_1[96]) );
  DFFRHQXL weight_1_reg_15__0_ ( .D(n14526), .CK(clk), .RN(rst_n), .Q(
        weight_1[90]) );
  DFFRHQXL weight_1_reg_14__0_ ( .D(n14525), .CK(clk), .RN(rst_n), .Q(
        weight_1[84]) );
  DFFRHQXL weight_1_reg_13__0_ ( .D(n14524), .CK(clk), .RN(rst_n), .Q(
        weight_1[78]) );
  DFFRHQXL weight_1_reg_12__0_ ( .D(n14523), .CK(clk), .RN(rst_n), .Q(
        weight_1[72]) );
  DFFRHQXL weight_1_reg_11__0_ ( .D(n14522), .CK(clk), .RN(rst_n), .Q(
        weight_1[66]) );
  DFFRHQXL weight_1_reg_10__0_ ( .D(n14521), .CK(clk), .RN(rst_n), .Q(
        weight_1[60]) );
  DFFRHQXL weight_1_reg_9__0_ ( .D(n14520), .CK(clk), .RN(rst_n), .Q(
        weight_1[54]) );
  DFFRHQXL weight_1_reg_8__0_ ( .D(n14519), .CK(clk), .RN(rst_n), .Q(
        weight_1[48]) );
  DFFRHQXL weight_1_reg_7__0_ ( .D(n14518), .CK(clk), .RN(rst_n), .Q(
        weight_1[42]) );
  DFFRHQXL weight_1_reg_6__0_ ( .D(n14517), .CK(clk), .RN(rst_n), .Q(
        weight_1[36]) );
  DFFRHQXL weight_1_reg_5__0_ ( .D(n14516), .CK(clk), .RN(rst_n), .Q(
        weight_1[30]) );
  DFFRHQXL weight_1_reg_4__0_ ( .D(n14515), .CK(clk), .RN(rst_n), .Q(
        weight_1[24]) );
  DFFRHQXL weight_1_reg_3__0_ ( .D(n14514), .CK(clk), .RN(rst_n), .Q(
        weight_1[18]) );
  DFFRHQXL weight_1_reg_2__0_ ( .D(n14513), .CK(clk), .RN(rst_n), .Q(
        weight_1[12]) );
  DFFRHQXL weight_1_reg_1__0_ ( .D(n14512), .CK(clk), .RN(rst_n), .Q(
        weight_1[6]) );
  DFFRHQXL weight_1_reg_0__0_ ( .D(n14511), .CK(clk), .RN(rst_n), .Q(
        weight_1[0]) );
  DFFRHQXL weight_1_reg_80__1_ ( .D(n14510), .CK(clk), .RN(rst_n), .Q(
        weight_1[481]) );
  DFFRHQXL weight_1_reg_79__1_ ( .D(n14509), .CK(clk), .RN(rst_n), .Q(
        weight_1[475]) );
  DFFRHQXL weight_1_reg_78__1_ ( .D(n14508), .CK(clk), .RN(rst_n), .Q(
        weight_1[469]) );
  DFFRHQXL weight_1_reg_77__1_ ( .D(n14507), .CK(clk), .RN(rst_n), .Q(
        weight_1[463]) );
  DFFRHQXL weight_1_reg_76__1_ ( .D(n14506), .CK(clk), .RN(rst_n), .Q(
        weight_1[457]) );
  DFFRHQXL weight_1_reg_75__1_ ( .D(n14505), .CK(clk), .RN(rst_n), .Q(
        weight_1[451]) );
  DFFRHQXL weight_1_reg_74__1_ ( .D(n14504), .CK(clk), .RN(rst_n), .Q(
        weight_1[445]) );
  DFFRHQXL weight_1_reg_73__1_ ( .D(n14503), .CK(clk), .RN(rst_n), .Q(
        weight_1[439]) );
  DFFRHQXL weight_1_reg_72__1_ ( .D(n14502), .CK(clk), .RN(rst_n), .Q(
        weight_1[433]) );
  DFFRHQXL weight_1_reg_71__1_ ( .D(n14501), .CK(clk), .RN(rst_n), .Q(
        weight_1[427]) );
  DFFRHQXL weight_1_reg_70__1_ ( .D(n14500), .CK(clk), .RN(rst_n), .Q(
        weight_1[421]) );
  DFFRHQXL weight_1_reg_69__1_ ( .D(n14499), .CK(clk), .RN(rst_n), .Q(
        weight_1[415]) );
  DFFRHQXL weight_1_reg_68__1_ ( .D(n14498), .CK(clk), .RN(rst_n), .Q(
        weight_1[409]) );
  DFFRHQXL weight_1_reg_67__1_ ( .D(n14497), .CK(clk), .RN(rst_n), .Q(
        weight_1[403]) );
  DFFRHQXL weight_1_reg_66__1_ ( .D(n14496), .CK(clk), .RN(rst_n), .Q(
        weight_1[397]) );
  DFFRHQXL weight_1_reg_65__1_ ( .D(n14495), .CK(clk), .RN(rst_n), .Q(
        weight_1[391]) );
  DFFRHQXL weight_1_reg_64__1_ ( .D(n14494), .CK(clk), .RN(rst_n), .Q(
        weight_1[385]) );
  DFFRHQXL weight_1_reg_63__1_ ( .D(n14493), .CK(clk), .RN(rst_n), .Q(
        weight_1[379]) );
  DFFRHQXL weight_1_reg_62__1_ ( .D(n14492), .CK(clk), .RN(rst_n), .Q(
        weight_1[373]) );
  DFFRHQXL weight_1_reg_61__1_ ( .D(n14491), .CK(clk), .RN(rst_n), .Q(
        weight_1[367]) );
  DFFRHQXL weight_1_reg_60__1_ ( .D(n14490), .CK(clk), .RN(rst_n), .Q(
        weight_1[361]) );
  DFFRHQXL weight_1_reg_59__1_ ( .D(n14489), .CK(clk), .RN(rst_n), .Q(
        weight_1[355]) );
  DFFRHQXL weight_1_reg_58__1_ ( .D(n14488), .CK(clk), .RN(rst_n), .Q(
        weight_1[349]) );
  DFFRHQXL weight_1_reg_57__1_ ( .D(n14487), .CK(clk), .RN(rst_n), .Q(
        weight_1[343]) );
  DFFRHQXL weight_1_reg_56__1_ ( .D(n14486), .CK(clk), .RN(rst_n), .Q(
        weight_1[337]) );
  DFFRHQXL weight_1_reg_55__1_ ( .D(n14485), .CK(clk), .RN(rst_n), .Q(
        weight_1[331]) );
  DFFRHQXL weight_1_reg_54__1_ ( .D(n14484), .CK(clk), .RN(rst_n), .Q(
        weight_1[325]) );
  DFFRHQXL weight_1_reg_53__1_ ( .D(n14483), .CK(clk), .RN(rst_n), .Q(
        weight_1[319]) );
  DFFRHQXL weight_1_reg_52__1_ ( .D(n14482), .CK(clk), .RN(rst_n), .Q(
        weight_1[313]) );
  DFFRHQXL weight_1_reg_51__1_ ( .D(n14481), .CK(clk), .RN(rst_n), .Q(
        weight_1[307]) );
  DFFRHQXL weight_1_reg_50__1_ ( .D(n14480), .CK(clk), .RN(rst_n), .Q(
        weight_1[301]) );
  DFFRHQXL weight_1_reg_49__1_ ( .D(n14479), .CK(clk), .RN(rst_n), .Q(
        weight_1[295]) );
  DFFRHQXL weight_1_reg_48__1_ ( .D(n14478), .CK(clk), .RN(rst_n), .Q(
        weight_1[289]) );
  DFFRHQXL weight_1_reg_47__1_ ( .D(n14477), .CK(clk), .RN(rst_n), .Q(
        weight_1[283]) );
  DFFRHQXL weight_1_reg_46__1_ ( .D(n14476), .CK(clk), .RN(rst_n), .Q(
        weight_1[277]) );
  DFFRHQXL weight_1_reg_45__1_ ( .D(n14475), .CK(clk), .RN(rst_n), .Q(
        weight_1[271]) );
  DFFRHQXL weight_1_reg_44__1_ ( .D(n14474), .CK(clk), .RN(rst_n), .Q(
        weight_1[265]) );
  DFFRHQXL weight_1_reg_43__1_ ( .D(n14473), .CK(clk), .RN(rst_n), .Q(
        weight_1[259]) );
  DFFRHQXL weight_1_reg_42__1_ ( .D(n14472), .CK(clk), .RN(rst_n), .Q(
        weight_1[253]) );
  DFFRHQXL weight_1_reg_41__1_ ( .D(n14471), .CK(clk), .RN(rst_n), .Q(
        weight_1[247]) );
  DFFRHQXL weight_1_reg_40__1_ ( .D(n14470), .CK(clk), .RN(rst_n), .Q(
        weight_1[241]) );
  DFFRHQXL weight_1_reg_39__1_ ( .D(n14469), .CK(clk), .RN(rst_n), .Q(
        weight_1[235]) );
  DFFRHQXL weight_1_reg_38__1_ ( .D(n14468), .CK(clk), .RN(rst_n), .Q(
        weight_1[229]) );
  DFFRHQXL weight_1_reg_37__1_ ( .D(n14467), .CK(clk), .RN(rst_n), .Q(
        weight_1[223]) );
  DFFRHQXL weight_1_reg_36__1_ ( .D(n14466), .CK(clk), .RN(rst_n), .Q(
        weight_1[217]) );
  DFFRHQXL weight_1_reg_35__1_ ( .D(n14465), .CK(clk), .RN(rst_n), .Q(
        weight_1[211]) );
  DFFRHQXL weight_1_reg_34__1_ ( .D(n14464), .CK(clk), .RN(rst_n), .Q(
        weight_1[205]) );
  DFFRHQXL weight_1_reg_33__1_ ( .D(n14463), .CK(clk), .RN(rst_n), .Q(
        weight_1[199]) );
  DFFRHQXL weight_1_reg_32__1_ ( .D(n14462), .CK(clk), .RN(rst_n), .Q(
        weight_1[193]) );
  DFFRHQXL weight_1_reg_31__1_ ( .D(n14461), .CK(clk), .RN(rst_n), .Q(
        weight_1[187]) );
  DFFRHQXL weight_1_reg_30__1_ ( .D(n14460), .CK(clk), .RN(rst_n), .Q(
        weight_1[181]) );
  DFFRHQXL weight_1_reg_29__1_ ( .D(n14459), .CK(clk), .RN(rst_n), .Q(
        weight_1[175]) );
  DFFRHQXL weight_1_reg_28__1_ ( .D(n14458), .CK(clk), .RN(rst_n), .Q(
        weight_1[169]) );
  DFFRHQXL weight_1_reg_27__1_ ( .D(n14457), .CK(clk), .RN(rst_n), .Q(
        weight_1[163]) );
  DFFRHQXL weight_1_reg_26__1_ ( .D(n14456), .CK(clk), .RN(rst_n), .Q(
        weight_1[157]) );
  DFFRHQXL weight_1_reg_25__1_ ( .D(n14455), .CK(clk), .RN(rst_n), .Q(
        weight_1[151]) );
  DFFRHQXL weight_1_reg_24__1_ ( .D(n14454), .CK(clk), .RN(rst_n), .Q(
        weight_1[145]) );
  DFFRHQXL weight_1_reg_23__1_ ( .D(n14453), .CK(clk), .RN(rst_n), .Q(
        weight_1[139]) );
  DFFRHQXL weight_1_reg_22__1_ ( .D(n14452), .CK(clk), .RN(rst_n), .Q(
        weight_1[133]) );
  DFFRHQXL weight_1_reg_21__1_ ( .D(n14451), .CK(clk), .RN(rst_n), .Q(
        weight_1[127]) );
  DFFRHQXL weight_1_reg_20__1_ ( .D(n14450), .CK(clk), .RN(rst_n), .Q(
        weight_1[121]) );
  DFFRHQXL weight_1_reg_19__1_ ( .D(n14449), .CK(clk), .RN(rst_n), .Q(
        weight_1[115]) );
  DFFRHQXL weight_1_reg_18__1_ ( .D(n14448), .CK(clk), .RN(rst_n), .Q(
        weight_1[109]) );
  DFFRHQXL weight_1_reg_17__1_ ( .D(n14447), .CK(clk), .RN(rst_n), .Q(
        weight_1[103]) );
  DFFRHQXL weight_1_reg_16__1_ ( .D(n14446), .CK(clk), .RN(rst_n), .Q(
        weight_1[97]) );
  DFFRHQXL weight_1_reg_15__1_ ( .D(n14445), .CK(clk), .RN(rst_n), .Q(
        weight_1[91]) );
  DFFRHQXL weight_1_reg_14__1_ ( .D(n14444), .CK(clk), .RN(rst_n), .Q(
        weight_1[85]) );
  DFFRHQXL weight_1_reg_13__1_ ( .D(n14443), .CK(clk), .RN(rst_n), .Q(
        weight_1[79]) );
  DFFRHQXL weight_1_reg_12__1_ ( .D(n14442), .CK(clk), .RN(rst_n), .Q(
        weight_1[73]) );
  DFFRHQXL weight_1_reg_11__1_ ( .D(n14441), .CK(clk), .RN(rst_n), .Q(
        weight_1[67]) );
  DFFRHQXL weight_1_reg_10__1_ ( .D(n14440), .CK(clk), .RN(rst_n), .Q(
        weight_1[61]) );
  DFFRHQXL weight_1_reg_9__1_ ( .D(n14439), .CK(clk), .RN(rst_n), .Q(
        weight_1[55]) );
  DFFRHQXL weight_1_reg_8__1_ ( .D(n14438), .CK(clk), .RN(rst_n), .Q(
        weight_1[49]) );
  DFFRHQXL weight_1_reg_7__1_ ( .D(n14437), .CK(clk), .RN(rst_n), .Q(
        weight_1[43]) );
  DFFRHQXL weight_1_reg_6__1_ ( .D(n14436), .CK(clk), .RN(rst_n), .Q(
        weight_1[37]) );
  DFFRHQXL weight_1_reg_5__1_ ( .D(n14435), .CK(clk), .RN(rst_n), .Q(
        weight_1[31]) );
  DFFRHQXL weight_1_reg_4__1_ ( .D(n14434), .CK(clk), .RN(rst_n), .Q(
        weight_1[25]) );
  DFFRHQXL weight_1_reg_3__1_ ( .D(n14433), .CK(clk), .RN(rst_n), .Q(
        weight_1[19]) );
  DFFRHQXL weight_1_reg_2__1_ ( .D(n14432), .CK(clk), .RN(rst_n), .Q(
        weight_1[13]) );
  DFFRHQXL weight_1_reg_1__1_ ( .D(n14431), .CK(clk), .RN(rst_n), .Q(
        weight_1[7]) );
  DFFRHQXL weight_1_reg_0__1_ ( .D(n14430), .CK(clk), .RN(rst_n), .Q(
        weight_1[1]) );
  DFFRHQXL weight_1_reg_80__2_ ( .D(n14429), .CK(clk), .RN(rst_n), .Q(
        weight_1[482]) );
  DFFRHQXL weight_1_reg_79__2_ ( .D(n14428), .CK(clk), .RN(rst_n), .Q(
        weight_1[476]) );
  DFFRHQXL weight_1_reg_78__2_ ( .D(n14427), .CK(clk), .RN(rst_n), .Q(
        weight_1[470]) );
  DFFRHQXL weight_1_reg_77__2_ ( .D(n14426), .CK(clk), .RN(rst_n), .Q(
        weight_1[464]) );
  DFFRHQXL weight_1_reg_76__2_ ( .D(n14425), .CK(clk), .RN(rst_n), .Q(
        weight_1[458]) );
  DFFRHQXL weight_1_reg_75__2_ ( .D(n14424), .CK(clk), .RN(rst_n), .Q(
        weight_1[452]) );
  DFFRHQXL weight_1_reg_74__2_ ( .D(n14423), .CK(clk), .RN(rst_n), .Q(
        weight_1[446]) );
  DFFRHQXL weight_1_reg_73__2_ ( .D(n14422), .CK(clk), .RN(rst_n), .Q(
        weight_1[440]) );
  DFFRHQXL weight_1_reg_72__2_ ( .D(n14421), .CK(clk), .RN(rst_n), .Q(
        weight_1[434]) );
  DFFRHQXL weight_1_reg_71__2_ ( .D(n14420), .CK(clk), .RN(rst_n), .Q(
        weight_1[428]) );
  DFFRHQXL weight_1_reg_70__2_ ( .D(n14419), .CK(clk), .RN(rst_n), .Q(
        weight_1[422]) );
  DFFRHQXL weight_1_reg_69__2_ ( .D(n14418), .CK(clk), .RN(rst_n), .Q(
        weight_1[416]) );
  DFFRHQXL weight_1_reg_68__2_ ( .D(n14417), .CK(clk), .RN(rst_n), .Q(
        weight_1[410]) );
  DFFRHQXL weight_1_reg_67__2_ ( .D(n14416), .CK(clk), .RN(rst_n), .Q(
        weight_1[404]) );
  DFFRHQXL weight_1_reg_66__2_ ( .D(n14415), .CK(clk), .RN(rst_n), .Q(
        weight_1[398]) );
  DFFRHQXL weight_1_reg_65__2_ ( .D(n14414), .CK(clk), .RN(rst_n), .Q(
        weight_1[392]) );
  DFFRHQXL weight_1_reg_64__2_ ( .D(n14413), .CK(clk), .RN(rst_n), .Q(
        weight_1[386]) );
  DFFRHQXL weight_1_reg_63__2_ ( .D(n14412), .CK(clk), .RN(rst_n), .Q(
        weight_1[380]) );
  DFFRHQXL weight_1_reg_62__2_ ( .D(n14411), .CK(clk), .RN(rst_n), .Q(
        weight_1[374]) );
  DFFRHQXL weight_1_reg_61__2_ ( .D(n14410), .CK(clk), .RN(rst_n), .Q(
        weight_1[368]) );
  DFFRHQXL weight_1_reg_60__2_ ( .D(n14409), .CK(clk), .RN(rst_n), .Q(
        weight_1[362]) );
  DFFRHQXL weight_1_reg_59__2_ ( .D(n14408), .CK(clk), .RN(rst_n), .Q(
        weight_1[356]) );
  DFFRHQXL weight_1_reg_58__2_ ( .D(n14407), .CK(clk), .RN(rst_n), .Q(
        weight_1[350]) );
  DFFRHQXL weight_1_reg_57__2_ ( .D(n14406), .CK(clk), .RN(rst_n), .Q(
        weight_1[344]) );
  DFFRHQXL weight_1_reg_56__2_ ( .D(n14405), .CK(clk), .RN(rst_n), .Q(
        weight_1[338]) );
  DFFRHQXL weight_1_reg_55__2_ ( .D(n14404), .CK(clk), .RN(rst_n), .Q(
        weight_1[332]) );
  DFFRHQXL weight_1_reg_54__2_ ( .D(n14403), .CK(clk), .RN(rst_n), .Q(
        weight_1[326]) );
  DFFRHQXL weight_1_reg_53__2_ ( .D(n14402), .CK(clk), .RN(rst_n), .Q(
        weight_1[320]) );
  DFFRHQXL weight_1_reg_52__2_ ( .D(n14401), .CK(clk), .RN(rst_n), .Q(
        weight_1[314]) );
  DFFRHQXL weight_1_reg_51__2_ ( .D(n14400), .CK(clk), .RN(rst_n), .Q(
        weight_1[308]) );
  DFFRHQXL weight_1_reg_50__2_ ( .D(n14399), .CK(clk), .RN(rst_n), .Q(
        weight_1[302]) );
  DFFRHQXL weight_1_reg_49__2_ ( .D(n14398), .CK(clk), .RN(rst_n), .Q(
        weight_1[296]) );
  DFFRHQXL weight_1_reg_48__2_ ( .D(n14397), .CK(clk), .RN(rst_n), .Q(
        weight_1[290]) );
  DFFRHQXL weight_1_reg_47__2_ ( .D(n14396), .CK(clk), .RN(rst_n), .Q(
        weight_1[284]) );
  DFFRHQXL weight_1_reg_46__2_ ( .D(n14395), .CK(clk), .RN(rst_n), .Q(
        weight_1[278]) );
  DFFRHQXL weight_1_reg_45__2_ ( .D(n14394), .CK(clk), .RN(rst_n), .Q(
        weight_1[272]) );
  DFFRHQXL weight_1_reg_44__2_ ( .D(n14393), .CK(clk), .RN(rst_n), .Q(
        weight_1[266]) );
  DFFRHQXL weight_1_reg_43__2_ ( .D(n14392), .CK(clk), .RN(rst_n), .Q(
        weight_1[260]) );
  DFFRHQXL weight_1_reg_42__2_ ( .D(n14391), .CK(clk), .RN(rst_n), .Q(
        weight_1[254]) );
  DFFRHQXL weight_1_reg_41__2_ ( .D(n14390), .CK(clk), .RN(rst_n), .Q(
        weight_1[248]) );
  DFFRHQXL weight_1_reg_40__2_ ( .D(n14389), .CK(clk), .RN(rst_n), .Q(
        weight_1[242]) );
  DFFRHQXL weight_1_reg_39__2_ ( .D(n14388), .CK(clk), .RN(rst_n), .Q(
        weight_1[236]) );
  DFFRHQXL weight_1_reg_38__2_ ( .D(n14387), .CK(clk), .RN(rst_n), .Q(
        weight_1[230]) );
  DFFRHQXL weight_1_reg_37__2_ ( .D(n14386), .CK(clk), .RN(rst_n), .Q(
        weight_1[224]) );
  DFFRHQXL weight_1_reg_36__2_ ( .D(n14385), .CK(clk), .RN(rst_n), .Q(
        weight_1[218]) );
  DFFRHQXL weight_1_reg_35__2_ ( .D(n14384), .CK(clk), .RN(rst_n), .Q(
        weight_1[212]) );
  DFFRHQXL weight_1_reg_34__2_ ( .D(n14383), .CK(clk), .RN(rst_n), .Q(
        weight_1[206]) );
  DFFRHQXL weight_1_reg_33__2_ ( .D(n14382), .CK(clk), .RN(rst_n), .Q(
        weight_1[200]) );
  DFFRHQXL weight_1_reg_32__2_ ( .D(n14381), .CK(clk), .RN(rst_n), .Q(
        weight_1[194]) );
  DFFRHQXL weight_1_reg_31__2_ ( .D(n14380), .CK(clk), .RN(rst_n), .Q(
        weight_1[188]) );
  DFFRHQXL weight_1_reg_30__2_ ( .D(n14379), .CK(clk), .RN(rst_n), .Q(
        weight_1[182]) );
  DFFRHQXL weight_1_reg_29__2_ ( .D(n14378), .CK(clk), .RN(rst_n), .Q(
        weight_1[176]) );
  DFFRHQXL weight_1_reg_28__2_ ( .D(n14377), .CK(clk), .RN(rst_n), .Q(
        weight_1[170]) );
  DFFRHQXL weight_1_reg_27__2_ ( .D(n14376), .CK(clk), .RN(rst_n), .Q(
        weight_1[164]) );
  DFFRHQXL weight_1_reg_26__2_ ( .D(n14375), .CK(clk), .RN(rst_n), .Q(
        weight_1[158]) );
  DFFRHQXL weight_1_reg_25__2_ ( .D(n14374), .CK(clk), .RN(rst_n), .Q(
        weight_1[152]) );
  DFFRHQXL weight_1_reg_24__2_ ( .D(n14373), .CK(clk), .RN(rst_n), .Q(
        weight_1[146]) );
  DFFRHQXL weight_1_reg_23__2_ ( .D(n14372), .CK(clk), .RN(rst_n), .Q(
        weight_1[140]) );
  DFFRHQXL weight_1_reg_22__2_ ( .D(n14371), .CK(clk), .RN(rst_n), .Q(
        weight_1[134]) );
  DFFRHQXL weight_1_reg_21__2_ ( .D(n14370), .CK(clk), .RN(rst_n), .Q(
        weight_1[128]) );
  DFFRHQXL weight_1_reg_20__2_ ( .D(n14369), .CK(clk), .RN(rst_n), .Q(
        weight_1[122]) );
  DFFRHQXL weight_1_reg_19__2_ ( .D(n14368), .CK(clk), .RN(rst_n), .Q(
        weight_1[116]) );
  DFFRHQXL weight_1_reg_18__2_ ( .D(n14367), .CK(clk), .RN(rst_n), .Q(
        weight_1[110]) );
  DFFRHQXL weight_1_reg_17__2_ ( .D(n14366), .CK(clk), .RN(rst_n), .Q(
        weight_1[104]) );
  DFFRHQXL weight_1_reg_16__2_ ( .D(n14365), .CK(clk), .RN(rst_n), .Q(
        weight_1[98]) );
  DFFRHQXL weight_1_reg_15__2_ ( .D(n14364), .CK(clk), .RN(rst_n), .Q(
        weight_1[92]) );
  DFFRHQXL weight_1_reg_14__2_ ( .D(n14363), .CK(clk), .RN(rst_n), .Q(
        weight_1[86]) );
  DFFRHQXL weight_1_reg_13__2_ ( .D(n14362), .CK(clk), .RN(rst_n), .Q(
        weight_1[80]) );
  DFFRHQXL weight_1_reg_12__2_ ( .D(n14361), .CK(clk), .RN(rst_n), .Q(
        weight_1[74]) );
  DFFRHQXL weight_1_reg_11__2_ ( .D(n14360), .CK(clk), .RN(rst_n), .Q(
        weight_1[68]) );
  DFFRHQXL weight_1_reg_10__2_ ( .D(n14359), .CK(clk), .RN(rst_n), .Q(
        weight_1[62]) );
  DFFRHQXL weight_1_reg_9__2_ ( .D(n14358), .CK(clk), .RN(rst_n), .Q(
        weight_1[56]) );
  DFFRHQXL weight_1_reg_8__2_ ( .D(n14357), .CK(clk), .RN(rst_n), .Q(
        weight_1[50]) );
  DFFRHQXL weight_1_reg_7__2_ ( .D(n14356), .CK(clk), .RN(rst_n), .Q(
        weight_1[44]) );
  DFFRHQXL weight_1_reg_6__2_ ( .D(n14355), .CK(clk), .RN(rst_n), .Q(
        weight_1[38]) );
  DFFRHQXL weight_1_reg_5__2_ ( .D(n14354), .CK(clk), .RN(rst_n), .Q(
        weight_1[32]) );
  DFFRHQXL weight_1_reg_4__2_ ( .D(n14353), .CK(clk), .RN(rst_n), .Q(
        weight_1[26]) );
  DFFRHQXL weight_1_reg_3__2_ ( .D(n14352), .CK(clk), .RN(rst_n), .Q(
        weight_1[20]) );
  DFFRHQXL weight_1_reg_2__2_ ( .D(n14351), .CK(clk), .RN(rst_n), .Q(
        weight_1[14]) );
  DFFRHQXL weight_1_reg_1__2_ ( .D(n14350), .CK(clk), .RN(rst_n), .Q(
        weight_1[8]) );
  DFFRHQXL weight_1_reg_0__2_ ( .D(n14349), .CK(clk), .RN(rst_n), .Q(
        weight_1[2]) );
  DFFRHQXL weight_1_reg_80__3_ ( .D(n14348), .CK(clk), .RN(rst_n), .Q(
        weight_1[483]) );
  DFFRHQXL weight_1_reg_79__3_ ( .D(n14347), .CK(clk), .RN(rst_n), .Q(
        weight_1[477]) );
  DFFRHQXL weight_1_reg_78__3_ ( .D(n14346), .CK(clk), .RN(rst_n), .Q(
        weight_1[471]) );
  DFFRHQXL weight_1_reg_77__3_ ( .D(n14345), .CK(clk), .RN(rst_n), .Q(
        weight_1[465]) );
  DFFRHQXL weight_1_reg_76__3_ ( .D(n14344), .CK(clk), .RN(rst_n), .Q(
        weight_1[459]) );
  DFFRHQXL weight_1_reg_75__3_ ( .D(n14343), .CK(clk), .RN(rst_n), .Q(
        weight_1[453]) );
  DFFRHQXL weight_1_reg_74__3_ ( .D(n14342), .CK(clk), .RN(rst_n), .Q(
        weight_1[447]) );
  DFFRHQXL weight_1_reg_73__3_ ( .D(n14341), .CK(clk), .RN(rst_n), .Q(
        weight_1[441]) );
  DFFRHQXL weight_1_reg_72__3_ ( .D(n14340), .CK(clk), .RN(rst_n), .Q(
        weight_1[435]) );
  DFFRHQXL weight_1_reg_71__3_ ( .D(n14339), .CK(clk), .RN(rst_n), .Q(
        weight_1[429]) );
  DFFRHQXL weight_1_reg_70__3_ ( .D(n14338), .CK(clk), .RN(rst_n), .Q(
        weight_1[423]) );
  DFFRHQXL weight_1_reg_69__3_ ( .D(n14337), .CK(clk), .RN(rst_n), .Q(
        weight_1[417]) );
  DFFRHQXL weight_1_reg_68__3_ ( .D(n14336), .CK(clk), .RN(rst_n), .Q(
        weight_1[411]) );
  DFFRHQXL weight_1_reg_67__3_ ( .D(n14335), .CK(clk), .RN(rst_n), .Q(
        weight_1[405]) );
  DFFRHQXL weight_1_reg_66__3_ ( .D(n14334), .CK(clk), .RN(rst_n), .Q(
        weight_1[399]) );
  DFFRHQXL weight_1_reg_65__3_ ( .D(n14333), .CK(clk), .RN(rst_n), .Q(
        weight_1[393]) );
  DFFRHQXL weight_1_reg_64__3_ ( .D(n14332), .CK(clk), .RN(rst_n), .Q(
        weight_1[387]) );
  DFFRHQXL weight_1_reg_63__3_ ( .D(n14331), .CK(clk), .RN(rst_n), .Q(
        weight_1[381]) );
  DFFRHQXL weight_1_reg_62__3_ ( .D(n14330), .CK(clk), .RN(rst_n), .Q(
        weight_1[375]) );
  DFFRHQXL weight_1_reg_61__3_ ( .D(n14329), .CK(clk), .RN(rst_n), .Q(
        weight_1[369]) );
  DFFRHQXL weight_1_reg_60__3_ ( .D(n14328), .CK(clk), .RN(rst_n), .Q(
        weight_1[363]) );
  DFFRHQXL weight_1_reg_59__3_ ( .D(n14327), .CK(clk), .RN(rst_n), .Q(
        weight_1[357]) );
  DFFRHQXL weight_1_reg_58__3_ ( .D(n14326), .CK(clk), .RN(rst_n), .Q(
        weight_1[351]) );
  DFFRHQXL weight_1_reg_57__3_ ( .D(n14325), .CK(clk), .RN(rst_n), .Q(
        weight_1[345]) );
  DFFRHQXL weight_1_reg_56__3_ ( .D(n14324), .CK(clk), .RN(rst_n), .Q(
        weight_1[339]) );
  DFFRHQXL weight_1_reg_55__3_ ( .D(n14323), .CK(clk), .RN(rst_n), .Q(
        weight_1[333]) );
  DFFRHQXL weight_1_reg_54__3_ ( .D(n14322), .CK(clk), .RN(rst_n), .Q(
        weight_1[327]) );
  DFFRHQXL weight_1_reg_53__3_ ( .D(n14321), .CK(clk), .RN(rst_n), .Q(
        weight_1[321]) );
  DFFRHQXL weight_1_reg_52__3_ ( .D(n14320), .CK(clk), .RN(rst_n), .Q(
        weight_1[315]) );
  DFFRHQXL weight_1_reg_51__3_ ( .D(n14319), .CK(clk), .RN(rst_n), .Q(
        weight_1[309]) );
  DFFRHQXL weight_1_reg_50__3_ ( .D(n14318), .CK(clk), .RN(rst_n), .Q(
        weight_1[303]) );
  DFFRHQXL weight_1_reg_49__3_ ( .D(n14317), .CK(clk), .RN(rst_n), .Q(
        weight_1[297]) );
  DFFRHQXL weight_1_reg_48__3_ ( .D(n14316), .CK(clk), .RN(rst_n), .Q(
        weight_1[291]) );
  DFFRHQXL weight_1_reg_47__3_ ( .D(n14315), .CK(clk), .RN(rst_n), .Q(
        weight_1[285]) );
  DFFRHQXL weight_1_reg_46__3_ ( .D(n14314), .CK(clk), .RN(rst_n), .Q(
        weight_1[279]) );
  DFFRHQXL weight_1_reg_45__3_ ( .D(n14313), .CK(clk), .RN(rst_n), .Q(
        weight_1[273]) );
  DFFRHQXL weight_1_reg_44__3_ ( .D(n14312), .CK(clk), .RN(rst_n), .Q(
        weight_1[267]) );
  DFFRHQXL weight_1_reg_43__3_ ( .D(n14311), .CK(clk), .RN(rst_n), .Q(
        weight_1[261]) );
  DFFRHQXL weight_1_reg_42__3_ ( .D(n14310), .CK(clk), .RN(rst_n), .Q(
        weight_1[255]) );
  DFFRHQXL weight_1_reg_41__3_ ( .D(n14309), .CK(clk), .RN(rst_n), .Q(
        weight_1[249]) );
  DFFRHQXL weight_1_reg_40__3_ ( .D(n14308), .CK(clk), .RN(rst_n), .Q(
        weight_1[243]) );
  DFFRHQXL weight_1_reg_39__3_ ( .D(n14307), .CK(clk), .RN(rst_n), .Q(
        weight_1[237]) );
  DFFRHQXL weight_1_reg_38__3_ ( .D(n14306), .CK(clk), .RN(rst_n), .Q(
        weight_1[231]) );
  DFFRHQXL weight_1_reg_37__3_ ( .D(n14305), .CK(clk), .RN(rst_n), .Q(
        weight_1[225]) );
  DFFRHQXL weight_1_reg_36__3_ ( .D(n14304), .CK(clk), .RN(rst_n), .Q(
        weight_1[219]) );
  DFFRHQXL weight_1_reg_35__3_ ( .D(n14303), .CK(clk), .RN(rst_n), .Q(
        weight_1[213]) );
  DFFRHQXL weight_1_reg_34__3_ ( .D(n14302), .CK(clk), .RN(rst_n), .Q(
        weight_1[207]) );
  DFFRHQXL weight_1_reg_33__3_ ( .D(n14301), .CK(clk), .RN(rst_n), .Q(
        weight_1[201]) );
  DFFRHQXL weight_1_reg_32__3_ ( .D(n14300), .CK(clk), .RN(rst_n), .Q(
        weight_1[195]) );
  DFFRHQXL weight_1_reg_31__3_ ( .D(n14299), .CK(clk), .RN(rst_n), .Q(
        weight_1[189]) );
  DFFRHQXL weight_1_reg_30__3_ ( .D(n14298), .CK(clk), .RN(rst_n), .Q(
        weight_1[183]) );
  DFFRHQXL weight_1_reg_29__3_ ( .D(n14297), .CK(clk), .RN(rst_n), .Q(
        weight_1[177]) );
  DFFRHQXL weight_1_reg_28__3_ ( .D(n14296), .CK(clk), .RN(rst_n), .Q(
        weight_1[171]) );
  DFFRHQXL weight_1_reg_27__3_ ( .D(n14295), .CK(clk), .RN(rst_n), .Q(
        weight_1[165]) );
  DFFRHQXL weight_1_reg_26__3_ ( .D(n14294), .CK(clk), .RN(rst_n), .Q(
        weight_1[159]) );
  DFFRHQXL weight_1_reg_25__3_ ( .D(n14293), .CK(clk), .RN(rst_n), .Q(
        weight_1[153]) );
  DFFRHQXL weight_1_reg_24__3_ ( .D(n14292), .CK(clk), .RN(rst_n), .Q(
        weight_1[147]) );
  DFFRHQXL weight_1_reg_23__3_ ( .D(n14291), .CK(clk), .RN(rst_n), .Q(
        weight_1[141]) );
  DFFRHQXL weight_1_reg_22__3_ ( .D(n14290), .CK(clk), .RN(rst_n), .Q(
        weight_1[135]) );
  DFFRHQXL weight_1_reg_21__3_ ( .D(n14289), .CK(clk), .RN(rst_n), .Q(
        weight_1[129]) );
  DFFRHQXL weight_1_reg_20__3_ ( .D(n14288), .CK(clk), .RN(rst_n), .Q(
        weight_1[123]) );
  DFFRHQXL weight_1_reg_19__3_ ( .D(n14287), .CK(clk), .RN(rst_n), .Q(
        weight_1[117]) );
  DFFRHQXL weight_1_reg_18__3_ ( .D(n14286), .CK(clk), .RN(rst_n), .Q(
        weight_1[111]) );
  DFFRHQXL weight_1_reg_17__3_ ( .D(n14285), .CK(clk), .RN(rst_n), .Q(
        weight_1[105]) );
  DFFRHQXL weight_1_reg_16__3_ ( .D(n14284), .CK(clk), .RN(rst_n), .Q(
        weight_1[99]) );
  DFFRHQXL weight_1_reg_15__3_ ( .D(n14283), .CK(clk), .RN(rst_n), .Q(
        weight_1[93]) );
  DFFRHQXL weight_1_reg_14__3_ ( .D(n14282), .CK(clk), .RN(rst_n), .Q(
        weight_1[87]) );
  DFFRHQXL weight_1_reg_13__3_ ( .D(n14281), .CK(clk), .RN(rst_n), .Q(
        weight_1[81]) );
  DFFRHQXL weight_1_reg_12__3_ ( .D(n14280), .CK(clk), .RN(rst_n), .Q(
        weight_1[75]) );
  DFFRHQXL weight_1_reg_11__3_ ( .D(n14279), .CK(clk), .RN(rst_n), .Q(
        weight_1[69]) );
  DFFRHQXL weight_1_reg_10__3_ ( .D(n14278), .CK(clk), .RN(rst_n), .Q(
        weight_1[63]) );
  DFFRHQXL weight_1_reg_9__3_ ( .D(n14277), .CK(clk), .RN(rst_n), .Q(
        weight_1[57]) );
  DFFRHQXL weight_1_reg_8__3_ ( .D(n14276), .CK(clk), .RN(rst_n), .Q(
        weight_1[51]) );
  DFFRHQXL weight_1_reg_7__3_ ( .D(n14275), .CK(clk), .RN(rst_n), .Q(
        weight_1[45]) );
  DFFRHQXL weight_1_reg_6__3_ ( .D(n14274), .CK(clk), .RN(rst_n), .Q(
        weight_1[39]) );
  DFFRHQXL weight_1_reg_5__3_ ( .D(n14273), .CK(clk), .RN(rst_n), .Q(
        weight_1[33]) );
  DFFRHQXL weight_1_reg_4__3_ ( .D(n14272), .CK(clk), .RN(rst_n), .Q(
        weight_1[27]) );
  DFFRHQXL weight_1_reg_3__3_ ( .D(n14271), .CK(clk), .RN(rst_n), .Q(
        weight_1[21]) );
  DFFRHQXL weight_1_reg_2__3_ ( .D(n14270), .CK(clk), .RN(rst_n), .Q(
        weight_1[15]) );
  DFFRHQXL weight_1_reg_1__3_ ( .D(n14269), .CK(clk), .RN(rst_n), .Q(
        weight_1[9]) );
  DFFRHQXL weight_1_reg_0__3_ ( .D(n14268), .CK(clk), .RN(rst_n), .Q(
        weight_1[3]) );
  DFFRHQXL weight_1_reg_80__4_ ( .D(n14267), .CK(clk), .RN(rst_n), .Q(
        weight_1[484]) );
  DFFRHQXL weight_1_reg_79__4_ ( .D(n14266), .CK(clk), .RN(rst_n), .Q(
        weight_1[478]) );
  DFFRHQXL weight_1_reg_78__4_ ( .D(n14265), .CK(clk), .RN(rst_n), .Q(
        weight_1[472]) );
  DFFRHQXL weight_1_reg_77__4_ ( .D(n14264), .CK(clk), .RN(rst_n), .Q(
        weight_1[466]) );
  DFFRHQXL weight_1_reg_76__4_ ( .D(n14263), .CK(clk), .RN(rst_n), .Q(
        weight_1[460]) );
  DFFRHQXL weight_1_reg_75__4_ ( .D(n14262), .CK(clk), .RN(rst_n), .Q(
        weight_1[454]) );
  DFFRHQXL weight_1_reg_74__4_ ( .D(n14261), .CK(clk), .RN(rst_n), .Q(
        weight_1[448]) );
  DFFRHQXL weight_1_reg_73__4_ ( .D(n14260), .CK(clk), .RN(rst_n), .Q(
        weight_1[442]) );
  DFFRHQXL weight_1_reg_72__4_ ( .D(n14259), .CK(clk), .RN(rst_n), .Q(
        weight_1[436]) );
  DFFRHQXL weight_1_reg_71__4_ ( .D(n14258), .CK(clk), .RN(rst_n), .Q(
        weight_1[430]) );
  DFFRHQXL weight_1_reg_70__4_ ( .D(n14257), .CK(clk), .RN(rst_n), .Q(
        weight_1[424]) );
  DFFRHQXL weight_1_reg_69__4_ ( .D(n14256), .CK(clk), .RN(rst_n), .Q(
        weight_1[418]) );
  DFFRHQXL weight_1_reg_68__4_ ( .D(n14255), .CK(clk), .RN(rst_n), .Q(
        weight_1[412]) );
  DFFRHQXL weight_1_reg_67__4_ ( .D(n14254), .CK(clk), .RN(rst_n), .Q(
        weight_1[406]) );
  DFFRHQXL weight_1_reg_66__4_ ( .D(n14253), .CK(clk), .RN(rst_n), .Q(
        weight_1[400]) );
  DFFRHQXL weight_1_reg_65__4_ ( .D(n14252), .CK(clk), .RN(rst_n), .Q(
        weight_1[394]) );
  DFFRHQXL weight_1_reg_64__4_ ( .D(n14251), .CK(clk), .RN(rst_n), .Q(
        weight_1[388]) );
  DFFRHQXL weight_1_reg_63__4_ ( .D(n14250), .CK(clk), .RN(rst_n), .Q(
        weight_1[382]) );
  DFFRHQXL weight_1_reg_62__4_ ( .D(n14249), .CK(clk), .RN(rst_n), .Q(
        weight_1[376]) );
  DFFRHQXL weight_1_reg_61__4_ ( .D(n14248), .CK(clk), .RN(rst_n), .Q(
        weight_1[370]) );
  DFFRHQXL weight_1_reg_60__4_ ( .D(n14247), .CK(clk), .RN(rst_n), .Q(
        weight_1[364]) );
  DFFRHQXL weight_1_reg_59__4_ ( .D(n14246), .CK(clk), .RN(rst_n), .Q(
        weight_1[358]) );
  DFFRHQXL weight_1_reg_58__4_ ( .D(n14245), .CK(clk), .RN(rst_n), .Q(
        weight_1[352]) );
  DFFRHQXL weight_1_reg_57__4_ ( .D(n14244), .CK(clk), .RN(rst_n), .Q(
        weight_1[346]) );
  DFFRHQXL weight_1_reg_56__4_ ( .D(n14243), .CK(clk), .RN(rst_n), .Q(
        weight_1[340]) );
  DFFRHQXL weight_1_reg_55__4_ ( .D(n14242), .CK(clk), .RN(rst_n), .Q(
        weight_1[334]) );
  DFFRHQXL weight_1_reg_54__4_ ( .D(n14241), .CK(clk), .RN(rst_n), .Q(
        weight_1[328]) );
  DFFRHQXL weight_1_reg_53__4_ ( .D(n14240), .CK(clk), .RN(rst_n), .Q(
        weight_1[322]) );
  DFFRHQXL weight_1_reg_52__4_ ( .D(n14239), .CK(clk), .RN(rst_n), .Q(
        weight_1[316]) );
  DFFRHQXL weight_1_reg_51__4_ ( .D(n14238), .CK(clk), .RN(rst_n), .Q(
        weight_1[310]) );
  DFFRHQXL weight_1_reg_50__4_ ( .D(n14237), .CK(clk), .RN(rst_n), .Q(
        weight_1[304]) );
  DFFRHQXL weight_1_reg_49__4_ ( .D(n14236), .CK(clk), .RN(rst_n), .Q(
        weight_1[298]) );
  DFFRHQXL weight_1_reg_48__4_ ( .D(n14235), .CK(clk), .RN(rst_n), .Q(
        weight_1[292]) );
  DFFRHQXL weight_1_reg_47__4_ ( .D(n14234), .CK(clk), .RN(rst_n), .Q(
        weight_1[286]) );
  DFFRHQXL weight_1_reg_46__4_ ( .D(n14233), .CK(clk), .RN(rst_n), .Q(
        weight_1[280]) );
  DFFRHQXL weight_1_reg_45__4_ ( .D(n14232), .CK(clk), .RN(rst_n), .Q(
        weight_1[274]) );
  DFFRHQXL weight_1_reg_44__4_ ( .D(n14231), .CK(clk), .RN(rst_n), .Q(
        weight_1[268]) );
  DFFRHQXL weight_1_reg_43__4_ ( .D(n14230), .CK(clk), .RN(rst_n), .Q(
        weight_1[262]) );
  DFFRHQXL weight_1_reg_42__4_ ( .D(n14229), .CK(clk), .RN(rst_n), .Q(
        weight_1[256]) );
  DFFRHQXL weight_1_reg_41__4_ ( .D(n14228), .CK(clk), .RN(rst_n), .Q(
        weight_1[250]) );
  DFFRHQXL weight_1_reg_40__4_ ( .D(n14227), .CK(clk), .RN(rst_n), .Q(
        weight_1[244]) );
  DFFRHQXL weight_1_reg_39__4_ ( .D(n14226), .CK(clk), .RN(rst_n), .Q(
        weight_1[238]) );
  DFFRHQXL weight_1_reg_38__4_ ( .D(n14225), .CK(clk), .RN(rst_n), .Q(
        weight_1[232]) );
  DFFRHQXL weight_1_reg_37__4_ ( .D(n14224), .CK(clk), .RN(rst_n), .Q(
        weight_1[226]) );
  DFFRHQXL weight_1_reg_36__4_ ( .D(n14223), .CK(clk), .RN(rst_n), .Q(
        weight_1[220]) );
  DFFRHQXL weight_1_reg_35__4_ ( .D(n14222), .CK(clk), .RN(rst_n), .Q(
        weight_1[214]) );
  DFFRHQXL weight_1_reg_34__4_ ( .D(n14221), .CK(clk), .RN(rst_n), .Q(
        weight_1[208]) );
  DFFRHQXL weight_1_reg_33__4_ ( .D(n14220), .CK(clk), .RN(rst_n), .Q(
        weight_1[202]) );
  DFFRHQXL weight_1_reg_32__4_ ( .D(n14219), .CK(clk), .RN(rst_n), .Q(
        weight_1[196]) );
  DFFRHQXL weight_1_reg_31__4_ ( .D(n14218), .CK(clk), .RN(rst_n), .Q(
        weight_1[190]) );
  DFFRHQXL weight_1_reg_30__4_ ( .D(n14217), .CK(clk), .RN(rst_n), .Q(
        weight_1[184]) );
  DFFRHQXL weight_1_reg_29__4_ ( .D(n14216), .CK(clk), .RN(rst_n), .Q(
        weight_1[178]) );
  DFFRHQXL weight_1_reg_28__4_ ( .D(n14215), .CK(clk), .RN(rst_n), .Q(
        weight_1[172]) );
  DFFRHQXL weight_1_reg_27__4_ ( .D(n14214), .CK(clk), .RN(rst_n), .Q(
        weight_1[166]) );
  DFFRHQXL weight_1_reg_26__4_ ( .D(n14213), .CK(clk), .RN(rst_n), .Q(
        weight_1[160]) );
  DFFRHQXL weight_1_reg_25__4_ ( .D(n14212), .CK(clk), .RN(rst_n), .Q(
        weight_1[154]) );
  DFFRHQXL weight_1_reg_24__4_ ( .D(n14211), .CK(clk), .RN(rst_n), .Q(
        weight_1[148]) );
  DFFRHQXL weight_1_reg_23__4_ ( .D(n14210), .CK(clk), .RN(rst_n), .Q(
        weight_1[142]) );
  DFFRHQXL weight_1_reg_22__4_ ( .D(n14209), .CK(clk), .RN(rst_n), .Q(
        weight_1[136]) );
  DFFRHQXL weight_1_reg_21__4_ ( .D(n14208), .CK(clk), .RN(rst_n), .Q(
        weight_1[130]) );
  DFFRHQXL weight_1_reg_20__4_ ( .D(n14207), .CK(clk), .RN(rst_n), .Q(
        weight_1[124]) );
  DFFRHQXL weight_1_reg_19__4_ ( .D(n14206), .CK(clk), .RN(rst_n), .Q(
        weight_1[118]) );
  DFFRHQXL weight_1_reg_18__4_ ( .D(n14205), .CK(clk), .RN(rst_n), .Q(
        weight_1[112]) );
  DFFRHQXL weight_1_reg_17__4_ ( .D(n14204), .CK(clk), .RN(rst_n), .Q(
        weight_1[106]) );
  DFFRHQXL weight_1_reg_16__4_ ( .D(n14203), .CK(clk), .RN(rst_n), .Q(
        weight_1[100]) );
  DFFRHQXL weight_1_reg_15__4_ ( .D(n14202), .CK(clk), .RN(rst_n), .Q(
        weight_1[94]) );
  DFFRHQXL weight_1_reg_14__4_ ( .D(n14201), .CK(clk), .RN(rst_n), .Q(
        weight_1[88]) );
  DFFRHQXL weight_1_reg_13__4_ ( .D(n14200), .CK(clk), .RN(rst_n), .Q(
        weight_1[82]) );
  DFFRHQXL weight_1_reg_12__4_ ( .D(n14199), .CK(clk), .RN(rst_n), .Q(
        weight_1[76]) );
  DFFRHQXL weight_1_reg_11__4_ ( .D(n14198), .CK(clk), .RN(rst_n), .Q(
        weight_1[70]) );
  DFFRHQXL weight_1_reg_10__4_ ( .D(n14197), .CK(clk), .RN(rst_n), .Q(
        weight_1[64]) );
  DFFRHQXL weight_1_reg_9__4_ ( .D(n14196), .CK(clk), .RN(rst_n), .Q(
        weight_1[58]) );
  DFFRHQXL weight_1_reg_8__4_ ( .D(n14195), .CK(clk), .RN(rst_n), .Q(
        weight_1[52]) );
  DFFRHQXL weight_1_reg_7__4_ ( .D(n14194), .CK(clk), .RN(rst_n), .Q(
        weight_1[46]) );
  DFFRHQXL weight_1_reg_6__4_ ( .D(n14193), .CK(clk), .RN(rst_n), .Q(
        weight_1[40]) );
  DFFRHQXL weight_1_reg_5__4_ ( .D(n14192), .CK(clk), .RN(rst_n), .Q(
        weight_1[34]) );
  DFFRHQXL weight_1_reg_4__4_ ( .D(n14191), .CK(clk), .RN(rst_n), .Q(
        weight_1[28]) );
  DFFRHQXL weight_1_reg_3__4_ ( .D(n14190), .CK(clk), .RN(rst_n), .Q(
        weight_1[22]) );
  DFFRHQXL weight_1_reg_2__4_ ( .D(n14189), .CK(clk), .RN(rst_n), .Q(
        weight_1[16]) );
  DFFRHQXL weight_1_reg_1__4_ ( .D(n14188), .CK(clk), .RN(rst_n), .Q(
        weight_1[10]) );
  DFFRHQXL weight_1_reg_0__4_ ( .D(n14187), .CK(clk), .RN(rst_n), .Q(
        weight_1[4]) );
  DFFRHQXL weight_1_reg_80__5_ ( .D(n14186), .CK(clk), .RN(rst_n), .Q(
        weight_1[485]) );
  DFFRHQXL weight_1_reg_79__5_ ( .D(n14185), .CK(clk), .RN(rst_n), .Q(
        weight_1[479]) );
  DFFRHQXL weight_1_reg_78__5_ ( .D(n14184), .CK(clk), .RN(rst_n), .Q(
        weight_1[473]) );
  DFFRHQXL weight_1_reg_77__5_ ( .D(n14183), .CK(clk), .RN(rst_n), .Q(
        weight_1[467]) );
  DFFRHQXL weight_1_reg_76__5_ ( .D(n14182), .CK(clk), .RN(rst_n), .Q(
        weight_1[461]) );
  DFFRHQXL weight_1_reg_75__5_ ( .D(n14181), .CK(clk), .RN(rst_n), .Q(
        weight_1[455]) );
  DFFRHQXL weight_1_reg_74__5_ ( .D(n14180), .CK(clk), .RN(rst_n), .Q(
        weight_1[449]) );
  DFFRHQXL weight_1_reg_73__5_ ( .D(n14179), .CK(clk), .RN(rst_n), .Q(
        weight_1[443]) );
  DFFRHQXL weight_1_reg_72__5_ ( .D(n14178), .CK(clk), .RN(rst_n), .Q(
        weight_1[437]) );
  DFFRHQXL weight_1_reg_71__5_ ( .D(n14177), .CK(clk), .RN(rst_n), .Q(
        weight_1[431]) );
  DFFRHQXL weight_1_reg_70__5_ ( .D(n14176), .CK(clk), .RN(rst_n), .Q(
        weight_1[425]) );
  DFFRHQXL weight_1_reg_69__5_ ( .D(n14175), .CK(clk), .RN(rst_n), .Q(
        weight_1[419]) );
  DFFRHQXL weight_1_reg_68__5_ ( .D(n14174), .CK(clk), .RN(rst_n), .Q(
        weight_1[413]) );
  DFFRHQXL weight_1_reg_67__5_ ( .D(n14173), .CK(clk), .RN(rst_n), .Q(
        weight_1[407]) );
  DFFRHQXL weight_1_reg_66__5_ ( .D(n14172), .CK(clk), .RN(rst_n), .Q(
        weight_1[401]) );
  DFFRHQXL weight_1_reg_65__5_ ( .D(n14171), .CK(clk), .RN(rst_n), .Q(
        weight_1[395]) );
  DFFRHQXL weight_1_reg_64__5_ ( .D(n14170), .CK(clk), .RN(rst_n), .Q(
        weight_1[389]) );
  DFFRHQXL weight_1_reg_63__5_ ( .D(n14169), .CK(clk), .RN(rst_n), .Q(
        weight_1[383]) );
  DFFRHQXL weight_1_reg_62__5_ ( .D(n14168), .CK(clk), .RN(rst_n), .Q(
        weight_1[377]) );
  DFFRHQXL weight_1_reg_61__5_ ( .D(n14167), .CK(clk), .RN(rst_n), .Q(
        weight_1[371]) );
  DFFRHQXL weight_1_reg_60__5_ ( .D(n14166), .CK(clk), .RN(rst_n), .Q(
        weight_1[365]) );
  DFFRHQXL weight_1_reg_59__5_ ( .D(n14165), .CK(clk), .RN(rst_n), .Q(
        weight_1[359]) );
  DFFRHQXL weight_1_reg_58__5_ ( .D(n14164), .CK(clk), .RN(rst_n), .Q(
        weight_1[353]) );
  DFFRHQXL weight_1_reg_57__5_ ( .D(n14163), .CK(clk), .RN(rst_n), .Q(
        weight_1[347]) );
  DFFRHQXL weight_1_reg_56__5_ ( .D(n14162), .CK(clk), .RN(rst_n), .Q(
        weight_1[341]) );
  DFFRHQXL weight_1_reg_55__5_ ( .D(n14161), .CK(clk), .RN(rst_n), .Q(
        weight_1[335]) );
  DFFRHQXL weight_1_reg_54__5_ ( .D(n14160), .CK(clk), .RN(rst_n), .Q(
        weight_1[329]) );
  DFFRHQXL weight_1_reg_53__5_ ( .D(n14159), .CK(clk), .RN(rst_n), .Q(
        weight_1[323]) );
  DFFRHQXL weight_1_reg_52__5_ ( .D(n14158), .CK(clk), .RN(rst_n), .Q(
        weight_1[317]) );
  DFFRHQXL weight_1_reg_51__5_ ( .D(n14157), .CK(clk), .RN(rst_n), .Q(
        weight_1[311]) );
  DFFRHQXL weight_1_reg_50__5_ ( .D(n14156), .CK(clk), .RN(rst_n), .Q(
        weight_1[305]) );
  DFFRHQXL weight_1_reg_49__5_ ( .D(n14155), .CK(clk), .RN(rst_n), .Q(
        weight_1[299]) );
  DFFRHQXL weight_1_reg_48__5_ ( .D(n14154), .CK(clk), .RN(rst_n), .Q(
        weight_1[293]) );
  DFFRHQXL weight_1_reg_47__5_ ( .D(n14153), .CK(clk), .RN(rst_n), .Q(
        weight_1[287]) );
  DFFRHQXL weight_1_reg_46__5_ ( .D(n14152), .CK(clk), .RN(rst_n), .Q(
        weight_1[281]) );
  DFFRHQXL weight_1_reg_45__5_ ( .D(n14151), .CK(clk), .RN(rst_n), .Q(
        weight_1[275]) );
  DFFRHQXL weight_1_reg_44__5_ ( .D(n14150), .CK(clk), .RN(rst_n), .Q(
        weight_1[269]) );
  DFFRHQXL weight_1_reg_43__5_ ( .D(n14149), .CK(clk), .RN(rst_n), .Q(
        weight_1[263]) );
  DFFRHQXL weight_1_reg_42__5_ ( .D(n14148), .CK(clk), .RN(rst_n), .Q(
        weight_1[257]) );
  DFFRHQXL weight_1_reg_41__5_ ( .D(n14147), .CK(clk), .RN(rst_n), .Q(
        weight_1[251]) );
  DFFRHQXL weight_1_reg_40__5_ ( .D(n14146), .CK(clk), .RN(rst_n), .Q(
        weight_1[245]) );
  DFFRHQXL weight_1_reg_39__5_ ( .D(n14145), .CK(clk), .RN(rst_n), .Q(
        weight_1[239]) );
  DFFRHQXL weight_1_reg_38__5_ ( .D(n14144), .CK(clk), .RN(rst_n), .Q(
        weight_1[233]) );
  DFFRHQXL weight_1_reg_37__5_ ( .D(n14143), .CK(clk), .RN(rst_n), .Q(
        weight_1[227]) );
  DFFRHQXL weight_1_reg_36__5_ ( .D(n14142), .CK(clk), .RN(rst_n), .Q(
        weight_1[221]) );
  DFFRHQXL weight_1_reg_35__5_ ( .D(n14141), .CK(clk), .RN(rst_n), .Q(
        weight_1[215]) );
  DFFRHQXL weight_1_reg_34__5_ ( .D(n14140), .CK(clk), .RN(rst_n), .Q(
        weight_1[209]) );
  DFFRHQXL weight_1_reg_33__5_ ( .D(n14139), .CK(clk), .RN(rst_n), .Q(
        weight_1[203]) );
  DFFRHQXL weight_1_reg_32__5_ ( .D(n14138), .CK(clk), .RN(rst_n), .Q(
        weight_1[197]) );
  DFFRHQXL weight_1_reg_31__5_ ( .D(n14137), .CK(clk), .RN(rst_n), .Q(
        weight_1[191]) );
  DFFRHQXL weight_1_reg_30__5_ ( .D(n14136), .CK(clk), .RN(rst_n), .Q(
        weight_1[185]) );
  DFFRHQXL weight_1_reg_29__5_ ( .D(n14135), .CK(clk), .RN(rst_n), .Q(
        weight_1[179]) );
  DFFRHQXL weight_1_reg_28__5_ ( .D(n14134), .CK(clk), .RN(rst_n), .Q(
        weight_1[173]) );
  DFFRHQXL weight_1_reg_27__5_ ( .D(n14133), .CK(clk), .RN(rst_n), .Q(
        weight_1[167]) );
  DFFRHQXL weight_1_reg_26__5_ ( .D(n14132), .CK(clk), .RN(rst_n), .Q(
        weight_1[161]) );
  DFFRHQXL weight_1_reg_25__5_ ( .D(n14131), .CK(clk), .RN(rst_n), .Q(
        weight_1[155]) );
  DFFRHQXL weight_1_reg_24__5_ ( .D(n14130), .CK(clk), .RN(rst_n), .Q(
        weight_1[149]) );
  DFFRHQXL weight_1_reg_23__5_ ( .D(n14129), .CK(clk), .RN(rst_n), .Q(
        weight_1[143]) );
  DFFRHQXL weight_1_reg_22__5_ ( .D(n14128), .CK(clk), .RN(rst_n), .Q(
        weight_1[137]) );
  DFFRHQXL weight_1_reg_21__5_ ( .D(n14127), .CK(clk), .RN(rst_n), .Q(
        weight_1[131]) );
  DFFRHQXL weight_1_reg_20__5_ ( .D(n14126), .CK(clk), .RN(rst_n), .Q(
        weight_1[125]) );
  DFFRHQXL weight_1_reg_19__5_ ( .D(n14125), .CK(clk), .RN(rst_n), .Q(
        weight_1[119]) );
  DFFRHQXL weight_1_reg_18__5_ ( .D(n14124), .CK(clk), .RN(rst_n), .Q(
        weight_1[113]) );
  DFFRHQXL weight_1_reg_17__5_ ( .D(n14123), .CK(clk), .RN(rst_n), .Q(
        weight_1[107]) );
  DFFRHQXL weight_1_reg_16__5_ ( .D(n14122), .CK(clk), .RN(rst_n), .Q(
        weight_1[101]) );
  DFFRHQXL weight_1_reg_15__5_ ( .D(n14121), .CK(clk), .RN(rst_n), .Q(
        weight_1[95]) );
  DFFRHQXL weight_1_reg_14__5_ ( .D(n14120), .CK(clk), .RN(rst_n), .Q(
        weight_1[89]) );
  DFFRHQXL weight_1_reg_13__5_ ( .D(n14119), .CK(clk), .RN(rst_n), .Q(
        weight_1[83]) );
  DFFRHQXL weight_1_reg_12__5_ ( .D(n14118), .CK(clk), .RN(rst_n), .Q(
        weight_1[77]) );
  DFFRHQXL weight_1_reg_11__5_ ( .D(n14117), .CK(clk), .RN(rst_n), .Q(
        weight_1[71]) );
  DFFRHQXL weight_1_reg_10__5_ ( .D(n14116), .CK(clk), .RN(rst_n), .Q(
        weight_1[65]) );
  DFFRHQXL weight_1_reg_9__5_ ( .D(n14115), .CK(clk), .RN(rst_n), .Q(
        weight_1[59]) );
  DFFRHQXL weight_1_reg_8__5_ ( .D(n14114), .CK(clk), .RN(rst_n), .Q(
        weight_1[53]) );
  DFFRHQXL weight_1_reg_7__5_ ( .D(n14113), .CK(clk), .RN(rst_n), .Q(
        weight_1[47]) );
  DFFRHQXL weight_1_reg_6__5_ ( .D(n14112), .CK(clk), .RN(rst_n), .Q(
        weight_1[41]) );
  DFFRHQXL weight_1_reg_5__5_ ( .D(n14111), .CK(clk), .RN(rst_n), .Q(
        weight_1[35]) );
  DFFRHQXL weight_1_reg_4__5_ ( .D(n14110), .CK(clk), .RN(rst_n), .Q(
        weight_1[29]) );
  DFFRHQXL weight_1_reg_3__5_ ( .D(n14109), .CK(clk), .RN(rst_n), .Q(
        weight_1[23]) );
  DFFRHQXL weight_1_reg_2__5_ ( .D(n14108), .CK(clk), .RN(rst_n), .Q(
        weight_1[17]) );
  DFFRHQXL weight_1_reg_1__5_ ( .D(n14107), .CK(clk), .RN(rst_n), .Q(
        weight_1[11]) );
  DFFRHQXL weight_1_reg_0__5_ ( .D(n14106), .CK(clk), .RN(rst_n), .Q(
        weight_1[5]) );
  DFFRHQXL weight_1_bias_3_reg_0_ ( .D(n14105), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_3[0]) );
  DFFRHQXL weight_1_bias_2_reg_0_ ( .D(n14104), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_2[0]) );
  DFFRHQXL weight_1_bias_1_reg_0_ ( .D(n14103), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_1[0]) );
  DFFRHQXL weight_1_bias_3_reg_1_ ( .D(n14102), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_3[1]) );
  DFFRHQXL weight_1_bias_2_reg_1_ ( .D(n14101), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_2[1]) );
  DFFRHQXL weight_1_bias_1_reg_1_ ( .D(n14100), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_1[1]) );
  DFFRHQXL weight_1_bias_3_reg_2_ ( .D(n14099), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_3[2]) );
  DFFRHQXL weight_1_bias_2_reg_2_ ( .D(n14098), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_2[2]) );
  DFFRHQXL weight_1_bias_1_reg_2_ ( .D(n14097), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_1[2]) );
  DFFRHQXL weight_1_bias_3_reg_3_ ( .D(n14096), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_3[3]) );
  DFFRHQXL weight_1_bias_2_reg_3_ ( .D(n14095), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_2[3]) );
  DFFRHQXL weight_1_bias_1_reg_3_ ( .D(n14094), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_1[3]) );
  DFFRHQXL weight_1_bias_3_reg_4_ ( .D(n14093), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_3[4]) );
  DFFRHQXL weight_1_bias_2_reg_4_ ( .D(n14092), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_2[4]) );
  DFFRHQXL weight_1_bias_1_reg_4_ ( .D(n14091), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_1[4]) );
  DFFRHQXL weight_1_bias_3_reg_5_ ( .D(n14090), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_3[5]) );
  DFFRHQXL affine_1_reg_2__9_ ( .D(n16492), .CK(clk), .RN(rst_n), .Q(
        affine_1[29]) );
  DFFRHQXL affine_1_reg_2__0_ ( .D(n16501), .CK(clk), .RN(rst_n), .Q(
        affine_1[20]) );
  DFFRHQXL affine_1_reg_2__1_ ( .D(n16500), .CK(clk), .RN(rst_n), .Q(
        affine_1[21]) );
  DFFRHQXL affine_1_reg_2__2_ ( .D(n16499), .CK(clk), .RN(rst_n), .Q(
        affine_1[22]) );
  DFFRHQXL affine_1_reg_2__3_ ( .D(n16498), .CK(clk), .RN(rst_n), .Q(
        affine_1[23]) );
  DFFRHQXL affine_1_reg_2__4_ ( .D(n16497), .CK(clk), .RN(rst_n), .Q(
        affine_1[24]) );
  DFFRHQXL affine_1_reg_2__5_ ( .D(n16496), .CK(clk), .RN(rst_n), .Q(
        affine_1[25]) );
  DFFRHQXL affine_1_reg_2__6_ ( .D(n16495), .CK(clk), .RN(rst_n), .Q(
        affine_1[26]) );
  DFFRHQXL affine_1_reg_2__7_ ( .D(n16494), .CK(clk), .RN(rst_n), .Q(
        affine_1[27]) );
  DFFRHQXL affine_1_reg_2__8_ ( .D(n16493), .CK(clk), .RN(rst_n), .Q(
        affine_1[28]) );
  DFFRHQXL weight_1_bias_2_reg_5_ ( .D(n14089), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_2[5]) );
  DFFRHQXL affine_1_reg_1__9_ ( .D(n16482), .CK(clk), .RN(rst_n), .Q(
        affine_1[19]) );
  DFFRHQXL affine_1_reg_1__0_ ( .D(n16491), .CK(clk), .RN(rst_n), .Q(
        affine_1[10]) );
  DFFRHQXL affine_1_reg_1__1_ ( .D(n16490), .CK(clk), .RN(rst_n), .Q(
        affine_1[11]) );
  DFFRHQXL affine_1_reg_1__2_ ( .D(n16489), .CK(clk), .RN(rst_n), .Q(
        affine_1[12]) );
  DFFRHQXL affine_1_reg_1__3_ ( .D(n16488), .CK(clk), .RN(rst_n), .Q(
        affine_1[13]) );
  DFFRHQXL affine_1_reg_1__4_ ( .D(n16487), .CK(clk), .RN(rst_n), .Q(
        affine_1[14]) );
  DFFRHQXL affine_1_reg_1__5_ ( .D(n16486), .CK(clk), .RN(rst_n), .Q(
        affine_1[15]) );
  DFFRHQXL affine_1_reg_1__6_ ( .D(n16485), .CK(clk), .RN(rst_n), .Q(
        affine_1[16]) );
  DFFRHQXL affine_1_reg_1__7_ ( .D(n16484), .CK(clk), .RN(rst_n), .Q(
        affine_1[17]) );
  DFFRHQXL affine_1_reg_1__8_ ( .D(n16483), .CK(clk), .RN(rst_n), .Q(
        affine_1[18]) );
  DFFRHQXL weight_1_bias_1_reg_5_ ( .D(n14088), .CK(clk), .RN(rst_n), .Q(
        weight_1_bias_1[5]) );
  DFFRHQXL affine_1_reg_0__9_ ( .D(n16504), .CK(clk), .RN(rst_n), .Q(
        affine_1[9]) );
  DFFRHQXL affine_1_reg_0__0_ ( .D(n16513), .CK(clk), .RN(rst_n), .Q(
        affine_1[0]) );
  DFFRHQXL affine_1_reg_0__1_ ( .D(n16512), .CK(clk), .RN(rst_n), .Q(
        affine_1[1]) );
  DFFRHQXL affine_1_reg_0__2_ ( .D(n16511), .CK(clk), .RN(rst_n), .Q(
        affine_1[2]) );
  DFFRHQXL affine_1_reg_0__3_ ( .D(n16510), .CK(clk), .RN(rst_n), .Q(
        affine_1[3]) );
  DFFRHQXL affine_1_reg_0__4_ ( .D(n16509), .CK(clk), .RN(rst_n), .Q(
        affine_1[4]) );
  DFFRHQXL affine_1_reg_0__5_ ( .D(n16508), .CK(clk), .RN(rst_n), .Q(
        affine_1[5]) );
  DFFRHQXL affine_1_reg_0__6_ ( .D(n16507), .CK(clk), .RN(rst_n), .Q(
        affine_1[6]) );
  DFFRHQXL affine_1_reg_0__7_ ( .D(n16506), .CK(clk), .RN(rst_n), .Q(
        affine_1[7]) );
  DFFRHQXL affine_1_reg_0__8_ ( .D(n16505), .CK(clk), .RN(rst_n), .Q(
        affine_1[8]) );
  ADDHXL add_x_358_U6 ( .A(n36246), .B(n35269), .CO(add_x_358_n5), .S(N29496)
         );
  ADDFXL intadd_1_U2 ( .A(conv_1[425]), .B(intadd_1_B_2_), .CI(intadd_1_n2), 
        .CO(intadd_1_n1), .S(intadd_1_SUM_2_) );
  CMPR42X1 DP_OP_5171J1_127_4278_U38 ( .A(affine_2[4]), .B(
        DP_OP_5171J1_127_4278_n89), .C(DP_OP_5171J1_127_4278_n107), .D(
        DP_OP_5171J1_127_4278_n98), .ICI(DP_OP_5171J1_127_4278_n67), .S(
        DP_OP_5171J1_127_4278_n64), .ICO(DP_OP_5171J1_127_4278_n62), .CO(
        DP_OP_5171J1_127_4278_n63) );
  CMPR42X1 DP_OP_5171J1_127_4278_U36 ( .A(DP_OP_5171J1_127_4278_n97), .B(
        DP_OP_5171J1_127_4278_n76), .C(DP_OP_5171J1_127_4278_n88), .D(
        DP_OP_5171J1_127_4278_n61), .ICI(DP_OP_5171J1_127_4278_n62), .S(
        DP_OP_5171J1_127_4278_n59), .ICO(DP_OP_5171J1_127_4278_n57), .CO(
        DP_OP_5171J1_127_4278_n58) );
  CMPR42X1 DP_OP_5171J1_127_4278_U34 ( .A(DP_OP_5171J1_127_4278_n96), .B(
        DP_OP_5171J1_127_4278_n87), .C(DP_OP_5171J1_127_4278_n60), .D(
        DP_OP_5171J1_127_4278_n56), .ICI(DP_OP_5171J1_127_4278_n57), .S(
        DP_OP_5171J1_127_4278_n54), .ICO(DP_OP_5171J1_127_4278_n52), .CO(
        DP_OP_5171J1_127_4278_n53) );
  CMPR42X1 DP_OP_5171J1_127_4278_U32 ( .A(DP_OP_5171J1_127_4278_n95), .B(
        DP_OP_5171J1_127_4278_n86), .C(DP_OP_5171J1_127_4278_n55), .D(
        DP_OP_5171J1_127_4278_n51), .ICI(DP_OP_5171J1_127_4278_n52), .S(
        DP_OP_5171J1_127_4278_n49), .ICO(DP_OP_5171J1_127_4278_n47), .CO(
        DP_OP_5171J1_127_4278_n48) );
  CMPR42X1 DP_OP_5171J1_127_4278_U30 ( .A(DP_OP_5171J1_127_4278_n94), .B(
        DP_OP_5171J1_127_4278_n85), .C(DP_OP_5171J1_127_4278_n50), .D(
        DP_OP_5171J1_127_4278_n46), .ICI(DP_OP_5171J1_127_4278_n47), .S(
        DP_OP_5171J1_127_4278_n44), .ICO(DP_OP_5171J1_127_4278_n42), .CO(
        DP_OP_5171J1_127_4278_n43) );
  CMPR42X1 DP_OP_5171J1_127_4278_U28 ( .A(DP_OP_5171J1_127_4278_n93), .B(
        DP_OP_5171J1_127_4278_n84), .C(DP_OP_5171J1_127_4278_n45), .D(
        DP_OP_5171J1_127_4278_n41), .ICI(DP_OP_5171J1_127_4278_n42), .S(
        DP_OP_5171J1_127_4278_n39), .ICO(DP_OP_5171J1_127_4278_n37), .CO(
        DP_OP_5171J1_127_4278_n38) );
  CMPR42X1 DP_OP_5171J1_127_4278_U25 ( .A(DP_OP_5171J1_127_4278_n83), .B(
        DP_OP_5171J1_127_4278_n101), .C(DP_OP_5171J1_127_4278_n40), .D(
        DP_OP_5171J1_127_4278_n36), .ICI(DP_OP_5171J1_127_4278_n37), .S(
        DP_OP_5171J1_127_4278_n34), .ICO(DP_OP_5171J1_127_4278_n32), .CO(
        DP_OP_5171J1_127_4278_n33) );
  CMPR42X1 DP_OP_5171J1_127_4278_U23 ( .A(DP_OP_5171J1_127_4278_n31), .B(
        DP_OP_5171J1_127_4278_n91), .C(DP_OP_5171J1_127_4278_n82), .D(
        DP_OP_5171J1_127_4278_n35), .ICI(DP_OP_5171J1_127_4278_n32), .S(
        DP_OP_5171J1_127_4278_n29), .ICO(DP_OP_5171J1_127_4278_n27), .CO(
        DP_OP_5171J1_127_4278_n28) );
  CMPR42X1 DP_OP_5171J1_127_4278_U22 ( .A(affine_2[12]), .B(affine_2[11]), .C(
        DP_OP_5171J1_127_4278_n81), .D(DP_OP_5171J1_127_4278_n90), .ICI(
        DP_OP_5171J1_127_4278_n27), .S(DP_OP_5171J1_127_4278_n26), .ICO(
        DP_OP_5171J1_127_4278_n24), .CO(DP_OP_5171J1_127_4278_n25) );
  CMPR42X1 DP_OP_5170J1_126_4278_U36 ( .A(DP_OP_5170J1_126_4278_n97), .B(
        DP_OP_5170J1_126_4278_n76), .C(DP_OP_5170J1_126_4278_n88), .D(
        DP_OP_5170J1_126_4278_n61), .ICI(DP_OP_5170J1_126_4278_n62), .S(
        DP_OP_5170J1_126_4278_n59), .ICO(DP_OP_5170J1_126_4278_n57), .CO(
        DP_OP_5170J1_126_4278_n58) );
  CMPR42X1 DP_OP_5170J1_126_4278_U34 ( .A(DP_OP_5170J1_126_4278_n96), .B(
        DP_OP_5170J1_126_4278_n87), .C(DP_OP_5170J1_126_4278_n60), .D(
        DP_OP_5170J1_126_4278_n56), .ICI(DP_OP_5170J1_126_4278_n57), .S(
        DP_OP_5170J1_126_4278_n54), .ICO(DP_OP_5170J1_126_4278_n52), .CO(
        DP_OP_5170J1_126_4278_n53) );
  CMPR42X1 DP_OP_5170J1_126_4278_U32 ( .A(DP_OP_5170J1_126_4278_n95), .B(
        DP_OP_5170J1_126_4278_n86), .C(DP_OP_5170J1_126_4278_n55), .D(
        DP_OP_5170J1_126_4278_n51), .ICI(DP_OP_5170J1_126_4278_n52), .S(
        DP_OP_5170J1_126_4278_n49), .ICO(DP_OP_5170J1_126_4278_n47), .CO(
        DP_OP_5170J1_126_4278_n48) );
  CMPR42X1 DP_OP_5170J1_126_4278_U30 ( .A(DP_OP_5170J1_126_4278_n94), .B(
        DP_OP_5170J1_126_4278_n85), .C(DP_OP_5170J1_126_4278_n50), .D(
        DP_OP_5170J1_126_4278_n46), .ICI(DP_OP_5170J1_126_4278_n47), .S(
        DP_OP_5170J1_126_4278_n44), .ICO(DP_OP_5170J1_126_4278_n42), .CO(
        DP_OP_5170J1_126_4278_n43) );
  CMPR42X1 DP_OP_5170J1_126_4278_U28 ( .A(DP_OP_5170J1_126_4278_n93), .B(
        DP_OP_5170J1_126_4278_n84), .C(DP_OP_5170J1_126_4278_n45), .D(
        DP_OP_5170J1_126_4278_n41), .ICI(DP_OP_5170J1_126_4278_n42), .S(
        DP_OP_5170J1_126_4278_n39), .ICO(DP_OP_5170J1_126_4278_n37), .CO(
        DP_OP_5170J1_126_4278_n38) );
  CMPR42X1 DP_OP_5170J1_126_4278_U25 ( .A(DP_OP_5170J1_126_4278_n83), .B(
        DP_OP_5170J1_126_4278_n101), .C(DP_OP_5170J1_126_4278_n40), .D(
        DP_OP_5170J1_126_4278_n36), .ICI(DP_OP_5170J1_126_4278_n37), .S(
        DP_OP_5170J1_126_4278_n34), .ICO(DP_OP_5170J1_126_4278_n32), .CO(
        DP_OP_5170J1_126_4278_n33) );
  CMPR42X1 DP_OP_5170J1_126_4278_U23 ( .A(DP_OP_5170J1_126_4278_n31), .B(
        DP_OP_5170J1_126_4278_n91), .C(DP_OP_5170J1_126_4278_n82), .D(
        DP_OP_5170J1_126_4278_n35), .ICI(DP_OP_5170J1_126_4278_n32), .S(
        DP_OP_5170J1_126_4278_n29), .ICO(DP_OP_5170J1_126_4278_n27), .CO(
        DP_OP_5170J1_126_4278_n28) );
  CMPR42X1 DP_OP_5170J1_126_4278_U22 ( .A(affine_2[28]), .B(affine_2[27]), .C(
        DP_OP_5170J1_126_4278_n81), .D(DP_OP_5170J1_126_4278_n90), .ICI(
        DP_OP_5170J1_126_4278_n27), .S(DP_OP_5170J1_126_4278_n26), .ICO(
        DP_OP_5170J1_126_4278_n24), .CO(DP_OP_5170J1_126_4278_n25) );
  CMPR42X1 DP_OP_5169J1_125_4278_U38 ( .A(affine_2[36]), .B(
        DP_OP_5169J1_125_4278_n89), .C(DP_OP_5169J1_125_4278_n107), .D(
        DP_OP_5169J1_125_4278_n98), .ICI(DP_OP_5169J1_125_4278_n67), .S(
        DP_OP_5169J1_125_4278_n64), .ICO(DP_OP_5169J1_125_4278_n62), .CO(
        DP_OP_5169J1_125_4278_n63) );
  CMPR42X1 DP_OP_5169J1_125_4278_U36 ( .A(DP_OP_5169J1_125_4278_n97), .B(
        DP_OP_5169J1_125_4278_n76), .C(DP_OP_5169J1_125_4278_n88), .D(
        DP_OP_5169J1_125_4278_n61), .ICI(DP_OP_5169J1_125_4278_n62), .S(
        DP_OP_5169J1_125_4278_n59), .ICO(DP_OP_5169J1_125_4278_n57), .CO(
        DP_OP_5169J1_125_4278_n58) );
  CMPR42X1 DP_OP_5169J1_125_4278_U34 ( .A(DP_OP_5169J1_125_4278_n96), .B(
        DP_OP_5169J1_125_4278_n87), .C(DP_OP_5169J1_125_4278_n60), .D(
        DP_OP_5169J1_125_4278_n56), .ICI(DP_OP_5169J1_125_4278_n57), .S(
        DP_OP_5169J1_125_4278_n54), .ICO(DP_OP_5169J1_125_4278_n52), .CO(
        DP_OP_5169J1_125_4278_n53) );
  CMPR42X1 DP_OP_5169J1_125_4278_U32 ( .A(DP_OP_5169J1_125_4278_n95), .B(
        DP_OP_5169J1_125_4278_n86), .C(DP_OP_5169J1_125_4278_n55), .D(
        DP_OP_5169J1_125_4278_n51), .ICI(DP_OP_5169J1_125_4278_n52), .S(
        DP_OP_5169J1_125_4278_n49), .ICO(DP_OP_5169J1_125_4278_n47), .CO(
        DP_OP_5169J1_125_4278_n48) );
  CMPR42X1 DP_OP_5169J1_125_4278_U30 ( .A(DP_OP_5169J1_125_4278_n94), .B(
        DP_OP_5169J1_125_4278_n85), .C(DP_OP_5169J1_125_4278_n50), .D(
        DP_OP_5169J1_125_4278_n46), .ICI(DP_OP_5169J1_125_4278_n47), .S(
        DP_OP_5169J1_125_4278_n44), .ICO(DP_OP_5169J1_125_4278_n42), .CO(
        DP_OP_5169J1_125_4278_n43) );
  CMPR42X1 DP_OP_5169J1_125_4278_U28 ( .A(DP_OP_5169J1_125_4278_n93), .B(
        DP_OP_5169J1_125_4278_n84), .C(DP_OP_5169J1_125_4278_n45), .D(
        DP_OP_5169J1_125_4278_n41), .ICI(DP_OP_5169J1_125_4278_n42), .S(
        DP_OP_5169J1_125_4278_n39), .ICO(DP_OP_5169J1_125_4278_n37), .CO(
        DP_OP_5169J1_125_4278_n38) );
  CMPR42X1 DP_OP_5169J1_125_4278_U25 ( .A(DP_OP_5169J1_125_4278_n83), .B(
        DP_OP_5169J1_125_4278_n101), .C(DP_OP_5169J1_125_4278_n40), .D(
        DP_OP_5169J1_125_4278_n36), .ICI(DP_OP_5169J1_125_4278_n37), .S(
        DP_OP_5169J1_125_4278_n34), .ICO(DP_OP_5169J1_125_4278_n32), .CO(
        DP_OP_5169J1_125_4278_n33) );
  CMPR42X1 DP_OP_5169J1_125_4278_U23 ( .A(DP_OP_5169J1_125_4278_n31), .B(
        DP_OP_5169J1_125_4278_n91), .C(DP_OP_5169J1_125_4278_n82), .D(
        DP_OP_5169J1_125_4278_n35), .ICI(DP_OP_5169J1_125_4278_n32), .S(
        DP_OP_5169J1_125_4278_n29), .ICO(DP_OP_5169J1_125_4278_n27), .CO(
        DP_OP_5169J1_125_4278_n28) );
  CMPR42X1 DP_OP_5169J1_125_4278_U22 ( .A(affine_2[44]), .B(affine_2[43]), .C(
        DP_OP_5169J1_125_4278_n81), .D(DP_OP_5169J1_125_4278_n90), .ICI(
        DP_OP_5169J1_125_4278_n27), .S(DP_OP_5169J1_125_4278_n26), .ICO(
        DP_OP_5169J1_125_4278_n24), .CO(DP_OP_5169J1_125_4278_n25) );
  CMPR42X1 DP_OP_5168J1_124_9881_U25 ( .A(DP_OP_5168J1_124_9881_n78), .B(
        DP_OP_5168J1_124_9881_n63), .C(DP_OP_5168J1_124_9881_n73), .D(
        DP_OP_5168J1_124_9881_n48), .ICI(DP_OP_5168J1_124_9881_n45), .S(
        DP_OP_5168J1_124_9881_n43), .ICO(DP_OP_5168J1_124_9881_n41), .CO(
        DP_OP_5168J1_124_9881_n42) );
  CMPR42X1 DP_OP_5168J1_124_9881_U21 ( .A(DP_OP_5168J1_124_9881_n67), .B(
        DP_OP_5168J1_124_9881_n57), .C(DP_OP_5168J1_124_9881_n41), .D(
        DP_OP_5168J1_124_9881_n40), .ICI(DP_OP_5168J1_124_9881_n38), .S(
        DP_OP_5168J1_124_9881_n36), .ICO(DP_OP_5168J1_124_9881_n34), .CO(
        DP_OP_5168J1_124_9881_n35) );
  CMPR42X1 DP_OP_5168J1_124_9881_U19 ( .A(DP_OP_5168J1_124_9881_n33), .B(
        DP_OP_5168J1_124_9881_n66), .C(DP_OP_5168J1_124_9881_n61), .D(
        DP_OP_5168J1_124_9881_n56), .ICI(DP_OP_5168J1_124_9881_n39), .S(
        DP_OP_5168J1_124_9881_n31), .ICO(DP_OP_5168J1_124_9881_n29), .CO(
        DP_OP_5168J1_124_9881_n30) );
  CMPR42X1 DP_OP_5168J1_124_9881_U18 ( .A(DP_OP_5168J1_124_9881_n71), .B(
        DP_OP_5168J1_124_9881_n76), .C(DP_OP_5168J1_124_9881_n37), .D(
        DP_OP_5168J1_124_9881_n34), .ICI(DP_OP_5168J1_124_9881_n31), .S(
        DP_OP_5168J1_124_9881_n28), .ICO(DP_OP_5168J1_124_9881_n26), .CO(
        DP_OP_5168J1_124_9881_n27) );
  CMPR42X1 DP_OP_5168J1_124_9881_U17 ( .A(affine_1[5]), .B(affine_1[6]), .C(
        DP_OP_5168J1_124_9881_n60), .D(DP_OP_5168J1_124_9881_n70), .ICI(
        DP_OP_5168J1_124_9881_n29), .S(DP_OP_5168J1_124_9881_n25), .ICO(
        DP_OP_5168J1_124_9881_n23), .CO(DP_OP_5168J1_124_9881_n24) );
  CMPR42X1 DP_OP_5168J1_124_9881_U16 ( .A(DP_OP_5168J1_124_9881_n65), .B(
        DP_OP_5168J1_124_9881_n55), .C(DP_OP_5168J1_124_9881_n25), .D(
        DP_OP_5168J1_124_9881_n30), .ICI(DP_OP_5168J1_124_9881_n26), .S(
        DP_OP_5168J1_124_9881_n22), .ICO(DP_OP_5168J1_124_9881_n20), .CO(
        DP_OP_5168J1_124_9881_n21) );
  CMPR42X1 DP_OP_5168J1_124_9881_U14 ( .A(DP_OP_5168J1_124_9881_n54), .B(
        DP_OP_5168J1_124_9881_n23), .C(DP_OP_5168J1_124_9881_n19), .D(
        DP_OP_5168J1_124_9881_n24), .ICI(DP_OP_5168J1_124_9881_n20), .S(
        DP_OP_5168J1_124_9881_n17), .ICO(DP_OP_5168J1_124_9881_n15), .CO(
        DP_OP_5168J1_124_9881_n16) );
  CMPR42X1 DP_OP_5168J1_124_9881_U13 ( .A(affine_1[8]), .B(
        DP_OP_5168J1_124_9881_n58), .C(DP_OP_5168J1_124_9881_n53), .D(
        DP_OP_5168J1_124_9881_n18), .ICI(DP_OP_5168J1_124_9881_n15), .S(
        DP_OP_5168J1_124_9881_n14), .ICO(DP_OP_5168J1_124_9881_n12), .CO(
        DP_OP_5168J1_124_9881_n13) );
  CMPR42X1 DP_OP_5167J1_123_9881_U25 ( .A(DP_OP_5167J1_123_9881_n78), .B(
        DP_OP_5167J1_123_9881_n63), .C(DP_OP_5167J1_123_9881_n73), .D(
        DP_OP_5167J1_123_9881_n48), .ICI(DP_OP_5167J1_123_9881_n45), .S(
        DP_OP_5167J1_123_9881_n43), .ICO(DP_OP_5167J1_123_9881_n41), .CO(
        DP_OP_5167J1_123_9881_n42) );
  CMPR42X1 DP_OP_5167J1_123_9881_U21 ( .A(DP_OP_5167J1_123_9881_n67), .B(
        DP_OP_5167J1_123_9881_n57), .C(DP_OP_5167J1_123_9881_n41), .D(
        DP_OP_5167J1_123_9881_n40), .ICI(DP_OP_5167J1_123_9881_n38), .S(
        DP_OP_5167J1_123_9881_n36), .ICO(DP_OP_5167J1_123_9881_n34), .CO(
        DP_OP_5167J1_123_9881_n35) );
  CMPR42X1 DP_OP_5167J1_123_9881_U19 ( .A(DP_OP_5167J1_123_9881_n33), .B(
        DP_OP_5167J1_123_9881_n66), .C(DP_OP_5167J1_123_9881_n61), .D(
        DP_OP_5167J1_123_9881_n56), .ICI(DP_OP_5167J1_123_9881_n39), .S(
        DP_OP_5167J1_123_9881_n31), .ICO(DP_OP_5167J1_123_9881_n29), .CO(
        DP_OP_5167J1_123_9881_n30) );
  CMPR42X1 DP_OP_5167J1_123_9881_U18 ( .A(DP_OP_5167J1_123_9881_n71), .B(
        DP_OP_5167J1_123_9881_n76), .C(DP_OP_5167J1_123_9881_n37), .D(
        DP_OP_5167J1_123_9881_n34), .ICI(DP_OP_5167J1_123_9881_n31), .S(
        DP_OP_5167J1_123_9881_n28), .ICO(DP_OP_5167J1_123_9881_n26), .CO(
        DP_OP_5167J1_123_9881_n27) );
  CMPR42X1 DP_OP_5167J1_123_9881_U17 ( .A(affine_1[15]), .B(affine_1[16]), .C(
        DP_OP_5167J1_123_9881_n60), .D(DP_OP_5167J1_123_9881_n70), .ICI(
        DP_OP_5167J1_123_9881_n29), .S(DP_OP_5167J1_123_9881_n25), .ICO(
        DP_OP_5167J1_123_9881_n23), .CO(DP_OP_5167J1_123_9881_n24) );
  CMPR42X1 DP_OP_5167J1_123_9881_U16 ( .A(DP_OP_5167J1_123_9881_n65), .B(
        DP_OP_5167J1_123_9881_n55), .C(DP_OP_5167J1_123_9881_n25), .D(
        DP_OP_5167J1_123_9881_n30), .ICI(DP_OP_5167J1_123_9881_n26), .S(
        DP_OP_5167J1_123_9881_n22), .ICO(DP_OP_5167J1_123_9881_n20), .CO(
        DP_OP_5167J1_123_9881_n21) );
  CMPR42X1 DP_OP_5167J1_123_9881_U14 ( .A(DP_OP_5167J1_123_9881_n54), .B(
        DP_OP_5167J1_123_9881_n23), .C(DP_OP_5167J1_123_9881_n19), .D(
        DP_OP_5167J1_123_9881_n24), .ICI(DP_OP_5167J1_123_9881_n20), .S(
        DP_OP_5167J1_123_9881_n17), .ICO(DP_OP_5167J1_123_9881_n15), .CO(
        DP_OP_5167J1_123_9881_n16) );
  CMPR42X1 DP_OP_5167J1_123_9881_U13 ( .A(affine_1[18]), .B(
        DP_OP_5167J1_123_9881_n58), .C(DP_OP_5167J1_123_9881_n53), .D(
        DP_OP_5167J1_123_9881_n18), .ICI(DP_OP_5167J1_123_9881_n15), .S(
        DP_OP_5167J1_123_9881_n14), .ICO(DP_OP_5167J1_123_9881_n12), .CO(
        DP_OP_5167J1_123_9881_n13) );
  CMPR42X1 DP_OP_5166J1_122_9881_U25 ( .A(DP_OP_5166J1_122_9881_n78), .B(
        DP_OP_5166J1_122_9881_n63), .C(DP_OP_5166J1_122_9881_n73), .D(
        DP_OP_5166J1_122_9881_n48), .ICI(DP_OP_5166J1_122_9881_n45), .S(
        DP_OP_5166J1_122_9881_n43), .ICO(DP_OP_5166J1_122_9881_n41), .CO(
        DP_OP_5166J1_122_9881_n42) );
  CMPR42X1 DP_OP_5166J1_122_9881_U21 ( .A(DP_OP_5166J1_122_9881_n67), .B(
        DP_OP_5166J1_122_9881_n57), .C(DP_OP_5166J1_122_9881_n41), .D(
        DP_OP_5166J1_122_9881_n40), .ICI(DP_OP_5166J1_122_9881_n38), .S(
        DP_OP_5166J1_122_9881_n36), .ICO(DP_OP_5166J1_122_9881_n34), .CO(
        DP_OP_5166J1_122_9881_n35) );
  CMPR42X1 DP_OP_5166J1_122_9881_U19 ( .A(DP_OP_5166J1_122_9881_n33), .B(
        DP_OP_5166J1_122_9881_n66), .C(DP_OP_5166J1_122_9881_n61), .D(
        DP_OP_5166J1_122_9881_n56), .ICI(DP_OP_5166J1_122_9881_n39), .S(
        DP_OP_5166J1_122_9881_n31), .ICO(DP_OP_5166J1_122_9881_n29), .CO(
        DP_OP_5166J1_122_9881_n30) );
  CMPR42X1 DP_OP_5166J1_122_9881_U18 ( .A(DP_OP_5166J1_122_9881_n71), .B(
        DP_OP_5166J1_122_9881_n76), .C(DP_OP_5166J1_122_9881_n37), .D(
        DP_OP_5166J1_122_9881_n34), .ICI(DP_OP_5166J1_122_9881_n31), .S(
        DP_OP_5166J1_122_9881_n28), .ICO(DP_OP_5166J1_122_9881_n26), .CO(
        DP_OP_5166J1_122_9881_n27) );
  CMPR42X1 DP_OP_5166J1_122_9881_U17 ( .A(affine_1[25]), .B(affine_1[26]), .C(
        DP_OP_5166J1_122_9881_n60), .D(DP_OP_5166J1_122_9881_n70), .ICI(
        DP_OP_5166J1_122_9881_n29), .S(DP_OP_5166J1_122_9881_n25), .ICO(
        DP_OP_5166J1_122_9881_n23), .CO(DP_OP_5166J1_122_9881_n24) );
  CMPR42X1 DP_OP_5166J1_122_9881_U16 ( .A(DP_OP_5166J1_122_9881_n65), .B(
        DP_OP_5166J1_122_9881_n55), .C(DP_OP_5166J1_122_9881_n25), .D(
        DP_OP_5166J1_122_9881_n30), .ICI(DP_OP_5166J1_122_9881_n26), .S(
        DP_OP_5166J1_122_9881_n22), .ICO(DP_OP_5166J1_122_9881_n20), .CO(
        DP_OP_5166J1_122_9881_n21) );
  CMPR42X1 DP_OP_5166J1_122_9881_U14 ( .A(DP_OP_5166J1_122_9881_n54), .B(
        DP_OP_5166J1_122_9881_n23), .C(DP_OP_5166J1_122_9881_n19), .D(
        DP_OP_5166J1_122_9881_n24), .ICI(DP_OP_5166J1_122_9881_n20), .S(
        DP_OP_5166J1_122_9881_n17), .ICO(DP_OP_5166J1_122_9881_n15), .CO(
        DP_OP_5166J1_122_9881_n16) );
  CMPR42X1 DP_OP_5166J1_122_9881_U13 ( .A(affine_1[28]), .B(
        DP_OP_5166J1_122_9881_n58), .C(DP_OP_5166J1_122_9881_n53), .D(
        DP_OP_5166J1_122_9881_n18), .ICI(DP_OP_5166J1_122_9881_n15), .S(
        DP_OP_5166J1_122_9881_n14), .ICO(DP_OP_5166J1_122_9881_n12), .CO(
        DP_OP_5166J1_122_9881_n13) );
  DFFSX1 out_valid_reg ( .D(n36250), .CK(clk), .SN(rst_n), .QN(out_valid) );
  DFFSX1 counter_reg_0_ ( .D(n16636), .CK(clk), .SN(rst_n), .Q(counter[0]), 
        .QN(n36248) );
  DFFSX1 cs_reg_3_ ( .D(n36249), .CK(clk), .SN(rst_n), .Q(n36247), .QN(cs[3])
         );
  DFFRHQXL cursor_reg_5_ ( .D(n16643), .CK(clk), .RN(rst_n), .Q(cursor[5]) );
  DFFRHQXL number_6_reg ( .D(n14086), .CK(clk), .RN(rst_n), .Q(number_6) );
  ADDFXL intadd_2_U3 ( .A(conv_1[3]), .B(intadd_2_B_1_), .CI(intadd_2_n3), 
        .CO(intadd_2_n2), .S(intadd_2_SUM_1_) );
  DFFRHQX1 counter_reg_3_ ( .D(N30142), .CK(clk), .RN(rst_n), .Q(counter[3])
         );
  DFFRHQXL number_2_reg ( .D(n14087), .CK(clk), .RN(rst_n), .Q(number_2) );
  DFFRHQXL number_4_reg ( .D(n14085), .CK(clk), .RN(rst_n), .Q(number_4) );
  DFFRHQX2 cursor_reg_3_ ( .D(n16641), .CK(clk), .RN(rst_n), .Q(N18014) );
  ADDFXL intadd_1_U3 ( .A(conv_1[424]), .B(intadd_1_B_1_), .CI(intadd_1_n3), 
        .CO(intadd_1_n2), .S(intadd_1_SUM_1_) );
  ADDFXL intadd_0_U3 ( .A(conv_2[3]), .B(intadd_0_B_1_), .CI(intadd_0_n3), 
        .CO(intadd_0_n2), .S(intadd_0_SUM_1_) );
  ADDFXL intadd_1_U4 ( .A(conv_1[423]), .B(intadd_1_B_0_), .CI(intadd_1_CI), 
        .CO(intadd_1_n3), .S(intadd_1_SUM_0_) );
  ADDFXL intadd_0_U4 ( .A(conv_2[2]), .B(intadd_0_B_0_), .CI(intadd_0_CI), 
        .CO(intadd_0_n3), .S(intadd_0_SUM_0_) );
  ADDFXL intadd_2_U4 ( .A(conv_1[2]), .B(intadd_2_B_0_), .CI(intadd_2_CI), 
        .CO(intadd_2_n3), .S(intadd_2_SUM_0_) );
  ADDFXL intadd_0_U2 ( .A(conv_2[4]), .B(intadd_0_B_2_), .CI(intadd_0_n2), 
        .CO(intadd_0_n1), .S(intadd_0_SUM_2_) );
  ADDFXL intadd_2_U2 ( .A(conv_1[4]), .B(intadd_2_B_2_), .CI(intadd_2_n2), 
        .CO(intadd_2_n1), .S(intadd_2_SUM_2_) );
  DFFRHQX4 cursor_reg_1_ ( .D(n16639), .CK(clk), .RN(rst_n), .Q(N17708) );
  NOR2X1 U15463 ( .A(n35269), .B(n35268), .Y(n16638) );
  NOR2X1 U15464 ( .A(n36250), .B(n36240), .Y(n14086) );
  NOR2X1 U15465 ( .A(n35245), .B(n35244), .Y(n35246) );
  NOR2X1 U15466 ( .A(n34855), .B(n34854), .Y(n34856) );
  NOR2X1 U15467 ( .A(n35265), .B(n35256), .Y(n35268) );
  NOR2X1 U15468 ( .A(n34937), .B(n34936), .Y(n34938) );
  NOR2X1 U15469 ( .A(n23941), .B(n34389), .Y(n23942) );
  NOR2X1 U15470 ( .A(n23884), .B(n36009), .Y(n23885) );
  NOR2X1 U15471 ( .A(n30226), .B(n16654), .Y(n30215) );
  NOR2X1 U15472 ( .A(n30210), .B(n36001), .Y(n30211) );
  NOR2X1 U15473 ( .A(n29428), .B(n16658), .Y(n21107) );
  NOR2X1 U15474 ( .A(n27213), .B(n16658), .Y(n24939) );
  NOR2X1 U15475 ( .A(n24266), .B(n16658), .Y(n24267) );
  NOR2X1 U15476 ( .A(n26297), .B(n36042), .Y(n24539) );
  NOR2X1 U15477 ( .A(n33719), .B(n33718), .Y(n33715) );
  NOR2X1 U15478 ( .A(n33735), .B(n33734), .Y(n33731) );
  NOR2X1 U15479 ( .A(n33752), .B(n33726), .Y(n33723) );
  NOR2X1 U15480 ( .A(n33752), .B(n33751), .Y(n33748) );
  NOR2X1 U15481 ( .A(n33571), .B(n33570), .Y(n33567) );
  NOR2X1 U15482 ( .A(n24520), .B(n36001), .Y(n24521) );
  NOR2X1 U15483 ( .A(n23461), .B(n36001), .Y(n21795) );
  NOR2X1 U15484 ( .A(n23742), .B(n36001), .Y(n23743) );
  NOR2X1 U15485 ( .A(n23455), .B(n36042), .Y(n23456) );
  NOR2X1 U15486 ( .A(n24555), .B(n36042), .Y(n24556) );
  NOR2X1 U15487 ( .A(n25073), .B(n16655), .Y(n24675) );
  NOR2X1 U15488 ( .A(n24525), .B(n16654), .Y(n24526) );
  NOR2X1 U15489 ( .A(n24668), .B(n16654), .Y(n24669) );
  NOR2X1 U15490 ( .A(n34052), .B(n16654), .Y(n22868) );
  NOR2X1 U15491 ( .A(n16655), .B(n27473), .Y(n27475) );
  NOR2X1 U15492 ( .A(n24486), .B(n16655), .Y(n24487) );
  NOR2X1 U15493 ( .A(n20360), .B(n30350), .Y(n36114) );
  NOR2X1 U15494 ( .A(n23267), .B(n23266), .Y(n23269) );
  NOR2X1 U15495 ( .A(n23667), .B(n23666), .Y(n23669) );
  NOR2X1 U15496 ( .A(n30760), .B(n30759), .Y(n30762) );
  NOR2X1 U15497 ( .A(n24458), .B(n24459), .Y(n23263) );
  NOR2X1 U15498 ( .A(n34207), .B(n34205), .Y(n34204) );
  NOR2X1 U15499 ( .A(n34576), .B(n34574), .Y(n34573) );
  NOR2X1 U15500 ( .A(n24433), .B(n24432), .Y(n24435) );
  NOR2X1 U15501 ( .A(n30959), .B(n30956), .Y(n30955) );
  NOR2X1 U15502 ( .A(n31148), .B(n31147), .Y(n31150) );
  NOR2X1 U15503 ( .A(n29162), .B(n29161), .Y(n26156) );
  NOR2X1 U15504 ( .A(n31739), .B(n31738), .Y(n31741) );
  NOR2X1 U15505 ( .A(n26940), .B(n26939), .Y(n26942) );
  NOR2X1 U15506 ( .A(n23540), .B(n23539), .Y(n23542) );
  NOR2X1 U15507 ( .A(n27357), .B(n27356), .Y(n27359) );
  NOR2X1 U15508 ( .A(n29548), .B(n29547), .Y(n29550) );
  NOR2X1 U15509 ( .A(n31692), .B(n31693), .Y(n29686) );
  NOR2X1 U15510 ( .A(n29638), .B(n29637), .Y(n29640) );
  NOR2X1 U15511 ( .A(n26928), .B(n26927), .Y(n26930) );
  NOR2X1 U15512 ( .A(n27457), .B(n27456), .Y(n27459) );
  NOR2X1 U15513 ( .A(n29605), .B(n29606), .Y(n27856) );
  NOR2X1 U15514 ( .A(n31233), .B(n31232), .Y(n31235) );
  NOR2X1 U15515 ( .A(n30544), .B(n30543), .Y(n30546) );
  NOR2X1 U15516 ( .A(n28109), .B(n28108), .Y(n28111) );
  NOR2X1 U15517 ( .A(n30031), .B(n30030), .Y(n30033) );
  NOR2X1 U15518 ( .A(n23170), .B(n23169), .Y(n23172) );
  NOR2X1 U15519 ( .A(n26779), .B(n26778), .Y(n26517) );
  NOR2X1 U15520 ( .A(n27261), .B(n27260), .Y(n27263) );
  NOR2X1 U15521 ( .A(n27107), .B(n27106), .Y(n27109) );
  NOR2X1 U15522 ( .A(n27479), .B(n27478), .Y(n27481) );
  NOR2X1 U15523 ( .A(n33398), .B(n33401), .Y(n30675) );
  NOR2X1 U15524 ( .A(n23936), .B(n23935), .Y(n23938) );
  NOR2X1 U15525 ( .A(n29227), .B(n29228), .Y(n29199) );
  NOR2X1 U15526 ( .A(n30488), .B(n30487), .Y(n30490) );
  NOR2X1 U15527 ( .A(n31637), .B(n31636), .Y(n31639) );
  NOR2X1 U15528 ( .A(n29898), .B(n29897), .Y(n29900) );
  NOR2X1 U15529 ( .A(n22838), .B(n22837), .Y(n22840) );
  NOR2X1 U15530 ( .A(n28943), .B(n28942), .Y(n28945) );
  NOR2X1 U15531 ( .A(n29971), .B(n29973), .Y(n27222) );
  NOR2X1 U15532 ( .A(n30179), .B(n30178), .Y(n30181) );
  NOR2X1 U15533 ( .A(n31933), .B(n31932), .Y(n31929) );
  NOR2X1 U15534 ( .A(n34715), .B(n34714), .Y(n34716) );
  NOR2X1 U15535 ( .A(n23229), .B(n23573), .Y(n23231) );
  NOR2X1 U15536 ( .A(n30319), .B(n30318), .Y(n30321) );
  NOR2X1 U15537 ( .A(n29745), .B(n29746), .Y(n22185) );
  NOR2X1 U15538 ( .A(n29566), .B(n29565), .Y(n29568) );
  NOR2X1 U15539 ( .A(n29011), .B(n29010), .Y(n29013) );
  NOR2X1 U15540 ( .A(n32018), .B(n32019), .Y(n23635) );
  NOR2X1 U15541 ( .A(n32297), .B(n32296), .Y(n32299) );
  NOR2X1 U15542 ( .A(n28972), .B(n28971), .Y(n28974) );
  NOR2X1 U15543 ( .A(n29035), .B(n29034), .Y(n29037) );
  NOR2X1 U15544 ( .A(n28796), .B(n28797), .Y(n24028) );
  NOR2X1 U15545 ( .A(n27837), .B(n27836), .Y(n27839) );
  NOR2X1 U15546 ( .A(n29245), .B(n25264), .Y(n25263) );
  NOR2X1 U15547 ( .A(n28599), .B(n28600), .Y(n25440) );
  NOR2X1 U15548 ( .A(n34280), .B(n34278), .Y(n34277) );
  NOR2X1 U15549 ( .A(n34240), .B(n34239), .Y(n34242) );
  NOR2X1 U15550 ( .A(n34246), .B(n34245), .Y(n34248) );
  NOR2X1 U15551 ( .A(n34151), .B(n34150), .Y(n34153) );
  NOR2X1 U15552 ( .A(n24924), .B(n24922), .Y(n24921) );
  NOR2X1 U15553 ( .A(n30901), .B(n30900), .Y(n30903) );
  NOR2X1 U15554 ( .A(n33220), .B(n33221), .Y(n32040) );
  NOR2X1 U15555 ( .A(n34561), .B(n34559), .Y(n34558) );
  NOR2X1 U15556 ( .A(n32176), .B(n32177), .Y(n31219) );
  NOR2X1 U15557 ( .A(n29577), .B(n29578), .Y(n27749) );
  NOR2X1 U15558 ( .A(n29174), .B(n29173), .Y(n29176) );
  NOR2X1 U15559 ( .A(n31350), .B(n31349), .Y(n31352) );
  NOR2X1 U15560 ( .A(n31792), .B(n31791), .Y(n31794) );
  NOR2X1 U15561 ( .A(n29753), .B(n26136), .Y(n26135) );
  NOR2X1 U15562 ( .A(n29221), .B(n29222), .Y(n26324) );
  NOR2X1 U15563 ( .A(n33957), .B(n33955), .Y(n33954) );
  NOR2X1 U15564 ( .A(n30952), .B(n30950), .Y(n30949) );
  NOR2X1 U15565 ( .A(n29101), .B(n29100), .Y(n29103) );
  NOR2X1 U15566 ( .A(n29904), .B(n29903), .Y(n29906) );
  NOR2X1 U15567 ( .A(n31950), .B(n31949), .Y(n31952) );
  NOR2X1 U15568 ( .A(n34304), .B(n34302), .Y(n34301) );
  NOR2X1 U15569 ( .A(n28810), .B(n28809), .Y(n28812) );
  NOR2X1 U15570 ( .A(n27660), .B(n27661), .Y(n27657) );
  NOR2X1 U15571 ( .A(n28771), .B(n28769), .Y(n28768) );
  NOR2X1 U15572 ( .A(n27747), .B(n27745), .Y(n27743) );
  NOR2X1 U15573 ( .A(n31444), .B(n31443), .Y(n31446) );
  NOR2X1 U15574 ( .A(n29702), .B(n29701), .Y(n29704) );
  NOR2X1 U15575 ( .A(n23141), .B(n23140), .Y(n23143) );
  NOR2X1 U15576 ( .A(n27167), .B(n27166), .Y(n27169) );
  NOR2X1 U15577 ( .A(n29542), .B(n29541), .Y(n29544) );
  NOR2X1 U15578 ( .A(n28892), .B(n28893), .Y(n28135) );
  NOR2X1 U15579 ( .A(n29832), .B(n29833), .Y(n29007) );
  NOR2X1 U15580 ( .A(n32025), .B(n32026), .Y(n32022) );
  NOR2X1 U15581 ( .A(n27295), .B(n27294), .Y(n27297) );
  NOR2X1 U15582 ( .A(n28051), .B(n28050), .Y(n28053) );
  NOR2X1 U15583 ( .A(n33938), .B(n33936), .Y(n33935) );
  NOR2X1 U15584 ( .A(n34407), .B(n34405), .Y(n34404) );
  NOR2X1 U15585 ( .A(n34400), .B(n34398), .Y(n34397) );
  NOR2X1 U15586 ( .A(n30557), .B(n30556), .Y(n30559) );
  NOR2X1 U15587 ( .A(n30563), .B(n30562), .Y(n30565) );
  NOR2X1 U15588 ( .A(n30748), .B(n30747), .Y(n30750) );
  NOR2X1 U15589 ( .A(n30468), .B(n30467), .Y(n30470) );
  NOR2X1 U15590 ( .A(n29880), .B(n29879), .Y(n29882) );
  NOR2X1 U15591 ( .A(n29763), .B(n29762), .Y(n29765) );
  NOR2X1 U15592 ( .A(n33315), .B(n31063), .Y(n31062) );
  NOR2X1 U15593 ( .A(n31003), .B(n31002), .Y(n31005) );
  NOR2X1 U15594 ( .A(n26364), .B(n26363), .Y(n26366) );
  NOR2X1 U15595 ( .A(n30889), .B(n30888), .Y(n30891) );
  NOR2X1 U15596 ( .A(n30858), .B(n30857), .Y(n30860) );
  NOR2X1 U15597 ( .A(n34297), .B(n34294), .Y(n34293) );
  NOR2X1 U15598 ( .A(n30922), .B(n30920), .Y(n30919) );
  NOR2X1 U15599 ( .A(n34348), .B(n34346), .Y(n34345) );
  NOR2X1 U15600 ( .A(n26307), .B(n26305), .Y(n26304) );
  NOR2X1 U15601 ( .A(n34384), .B(n34381), .Y(n34380) );
  NOR2X1 U15602 ( .A(n27113), .B(n25239), .Y(n25238) );
  NOR2X1 U15603 ( .A(n27278), .B(intadd_2_n1), .Y(n27070) );
  NOR2X1 U15604 ( .A(n23923), .B(n26667), .Y(n23917) );
  NOR2X1 U15605 ( .A(n35732), .B(n33111), .Y(n31497) );
  NOR2X1 U15606 ( .A(n34529), .B(n34528), .Y(n34537) );
  NOR2X1 U15607 ( .A(n27386), .B(n27387), .Y(n27385) );
  NOR2X1 U15608 ( .A(n23998), .B(n23999), .Y(n23997) );
  NOR2X1 U15609 ( .A(n23867), .B(n23868), .Y(n23866) );
  NOR2X1 U15610 ( .A(n28965), .B(n28966), .Y(n28964) );
  NOR2X1 U15611 ( .A(n34570), .B(n34571), .Y(n29536) );
  NOR2X1 U15612 ( .A(n30191), .B(n29350), .Y(n29322) );
  NOR2X1 U15613 ( .A(n23492), .B(n23493), .Y(n23491) );
  NOR2X1 U15614 ( .A(n29935), .B(n31310), .Y(n29922) );
  NOR2X1 U15615 ( .A(n28644), .B(n24175), .Y(n24174) );
  NOR2X1 U15616 ( .A(n34132), .B(n34133), .Y(n33668) );
  NOR2X1 U15617 ( .A(n33842), .B(n31915), .Y(n31910) );
  NOR2X1 U15618 ( .A(n29364), .B(n29365), .Y(n29363) );
  NOR2X1 U15619 ( .A(n32557), .B(n32559), .Y(n19211) );
  NOR2X1 U15620 ( .A(n35339), .B(n26754), .Y(n19138) );
  NOR2X1 U15621 ( .A(n33780), .B(n31513), .Y(n19068) );
  NOR2X1 U15622 ( .A(n35463), .B(n33089), .Y(n19158) );
  NOR2X1 U15623 ( .A(n32887), .B(n29824), .Y(n18861) );
  NOR2X1 U15624 ( .A(n18997), .B(n30511), .Y(n30513) );
  NOR2X1 U15625 ( .A(n34823), .B(n25393), .Y(n25303) );
  NOR2X1 U15626 ( .A(n18997), .B(n30549), .Y(n30551) );
  NOR2X1 U15627 ( .A(conv_3[178]), .B(n32644), .Y(n32643) );
  NOR2X1 U15628 ( .A(n21944), .B(n24211), .Y(n21805) );
  NOR2X1 U15629 ( .A(n28191), .B(n28137), .Y(n19049) );
  NOR2X1 U15630 ( .A(n30536), .B(n30618), .Y(n30538) );
  NOR2X1 U15631 ( .A(n36088), .B(n27910), .Y(n18941) );
  NOR2X1 U15632 ( .A(n33979), .B(n28627), .Y(n19119) );
  NOR2X1 U15633 ( .A(n28644), .B(n28643), .Y(n28650) );
  NOR2X1 U15634 ( .A(n30940), .B(n30202), .Y(n19178) );
  NOR2X1 U15635 ( .A(ns[1]), .B(n19632), .Y(n20614) );
  NOR2X1 U15636 ( .A(n24040), .B(n22713), .Y(n20732) );
  AND4X2 U15637 ( .A(n26273), .B(n26272), .C(n26271), .D(n26288), .Y(n26287)
         );
  AND4X2 U15638 ( .A(n26655), .B(n26654), .C(n26653), .D(pool[19]), .Y(n26659)
         );
  AND4X2 U15639 ( .A(n21281), .B(n21280), .C(n21375), .D(n21374), .Y(n21379)
         );
  AND4X2 U15640 ( .A(n21782), .B(n21781), .C(n21780), .D(pool[24]), .Y(n21786)
         );
  NOR2X1 U15641 ( .A(conv_3[281]), .B(n31762), .Y(n32597) );
  AND4X2 U15642 ( .A(n28569), .B(n28568), .C(n28567), .D(n28589), .Y(n28588)
         );
  AND4X2 U15643 ( .A(n24796), .B(n24795), .C(n24794), .D(pool[64]), .Y(n24800)
         );
  NOR2X1 U15644 ( .A(n35639), .B(n31573), .Y(n35636) );
  AND4X2 U15645 ( .A(n24128), .B(n24119), .C(n24118), .D(n24117), .Y(n24127)
         );
  AND4X2 U15646 ( .A(n26483), .B(n26482), .C(n26481), .D(n26480), .Y(n26486)
         );
  NOR2X1 U15647 ( .A(conv_3[461]), .B(n31523), .Y(n31519) );
  NOR2X1 U15648 ( .A(conv_3[476]), .B(n32339), .Y(n32327) );
  AND4X2 U15649 ( .A(n25803), .B(n25794), .C(n25793), .D(n25792), .Y(n25801)
         );
  AND4X2 U15650 ( .A(n26106), .B(n26107), .C(n26101), .D(pool[84]), .Y(n26105)
         );
  AND4X2 U15651 ( .A(n20343), .B(n20331), .C(n20330), .D(n20329), .Y(n20342)
         );
  AND4X2 U15652 ( .A(n25195), .B(n25194), .C(n25193), .D(n25192), .Y(n25196)
         );
  AND4X2 U15653 ( .A(n21721), .B(n21720), .C(n21719), .D(n21718), .Y(n21722)
         );
  NOR2X1 U15654 ( .A(n18653), .B(n18652), .Y(n18721) );
  NOR2X1 U15655 ( .A(n30927), .B(n31002), .Y(n30925) );
  NOR2X1 U15656 ( .A(n31994), .B(n32010), .Y(n31998) );
  NOR2X1 U15657 ( .A(n28174), .B(n28176), .Y(n28172) );
  NOR2X1 U15658 ( .A(n31780), .B(n31779), .Y(n34195) );
  ADDFX2 U15659 ( .A(conv_3[132]), .B(n35622), .CI(n34757), .CO(n34784), .S(
        n33711) );
  NOR2X1 U15660 ( .A(conv_1[431]), .B(n35507), .Y(n29330) );
  NOR2X1 U15661 ( .A(conv_2[251]), .B(n35940), .Y(n29456) );
  NOR2X1 U15662 ( .A(conv_2[41]), .B(n29618), .Y(n27724) );
  NOR2X1 U15663 ( .A(conv_1[401]), .B(n35476), .Y(n35480) );
  NOR2X1 U15664 ( .A(conv_3[57]), .B(n33820), .Y(n33821) );
  NOR2X1 U15665 ( .A(conv_3[357]), .B(n33724), .Y(n33725) );
  NOR2X1 U15666 ( .A(conv_1[252]), .B(n33660), .Y(n33661) );
  NOR2X1 U15667 ( .A(conv_1[492]), .B(n30326), .Y(n33210) );
  NOR2X1 U15668 ( .A(n20168), .B(n20167), .Y(n20179) );
  AND4X2 U15669 ( .A(n25444), .B(n25024), .C(n25023), .D(n25022), .Y(n25025)
         );
  NOR2X1 U15670 ( .A(n35138), .B(n35137), .Y(n35251) );
  NOR2X1 U15671 ( .A(counter[5]), .B(n18773), .Y(n26848) );
  AND4X2 U15672 ( .A(n18425), .B(n18424), .C(n18423), .D(n18444), .Y(n18443)
         );
  AND4X2 U15673 ( .A(n25476), .B(n25475), .C(n25474), .D(n25473), .Y(n27369)
         );
  NOR2X1 U15674 ( .A(n25820), .B(n35196), .Y(n21978) );
  NOR2X1 U15675 ( .A(n21724), .B(n28575), .Y(n19775) );
  AND4X2 U15676 ( .A(n27980), .B(n26603), .C(n26602), .D(n26601), .Y(n26628)
         );
  INVX2 U15677 ( .A(ns[0]), .Y(n19242) );
  NOR2X1 U15678 ( .A(n25814), .B(n26474), .Y(n25818) );
  NOR2X1 U15679 ( .A(n25194), .B(n25193), .Y(n25191) );
  NOR2X1 U15680 ( .A(n35999), .B(n35994), .Y(n29611) );
  NOR2X1 U15681 ( .A(n21281), .B(n21280), .Y(n21377) );
  NOR2X1 U15682 ( .A(n20064), .B(n20063), .Y(n20093) );
  NOR2X1 U15683 ( .A(n26545), .B(n26544), .Y(n27978) );
  NOR2X1 U15684 ( .A(n28587), .B(n28569), .Y(n28542) );
  NOR2X1 U15685 ( .A(conv_2[191]), .B(n29904), .Y(n30948) );
  NOR2X1 U15686 ( .A(conv_1[71]), .B(n27089), .Y(n26311) );
  NOR2X1 U15687 ( .A(n21781), .B(n21782), .Y(n21699) );
  NOR2X1 U15688 ( .A(n25064), .B(n25063), .Y(n35364) );
  NOR2X1 U15689 ( .A(n31579), .B(n32221), .Y(n32222) );
  NOR2X1 U15690 ( .A(n21390), .B(n35198), .Y(n19530) );
  NOR2X1 U15691 ( .A(n23181), .B(n23186), .Y(n23188) );
  NOR2X1 U15692 ( .A(n29223), .B(n29328), .Y(n35507) );
  NOR2X1 U15693 ( .A(conv_1[221]), .B(n28599), .Y(n28601) );
  NOR2X1 U15694 ( .A(n26755), .B(n32780), .Y(n32784) );
  NOR2X1 U15695 ( .A(n33169), .B(n36081), .Y(n33172) );
  NOR2X1 U15696 ( .A(n25794), .B(n25793), .Y(n25778) );
  NOR2X1 U15697 ( .A(n29481), .B(n29480), .Y(n28120) );
  NOR2X1 U15698 ( .A(n28795), .B(n28791), .Y(n27921) );
  NOR2X1 U15699 ( .A(n35777), .B(n35774), .Y(n31725) );
  NOR2X1 U15700 ( .A(n35617), .B(n35614), .Y(n32114) );
  NOR2X1 U15701 ( .A(n35609), .B(n35606), .Y(n31817) );
  NOR2X1 U15702 ( .A(n32081), .B(n32077), .Y(n32346) );
  NOR2X1 U15703 ( .A(n36083), .B(n36080), .Y(n36087) );
  NOR2X1 U15704 ( .A(n33464), .B(n32789), .Y(n33967) );
  NOR2X1 U15705 ( .A(n29119), .B(n35700), .Y(n35705) );
  NOR2X1 U15706 ( .A(n30243), .B(n30242), .Y(n33732) );
  NOR2X1 U15707 ( .A(n24891), .B(n24904), .Y(n24894) );
  NOR2X1 U15708 ( .A(n27160), .B(n27165), .Y(n35514) );
  NOR2X1 U15709 ( .A(n24729), .B(n24728), .Y(n26150) );
  NOR2X1 U15710 ( .A(n35441), .B(n35442), .Y(n35440) );
  NOR2X1 U15711 ( .A(n35111), .B(n35110), .Y(n35253) );
  NOR2X1 U15712 ( .A(n26578), .B(n26577), .Y(n27980) );
  NOR2X1 U15713 ( .A(n20752), .B(n20751), .Y(n25822) );
  NOR2X1 U15714 ( .A(n30214), .B(n30212), .Y(n30210) );
  NOR2X1 U15715 ( .A(n27239), .B(n30030), .Y(n30043) );
  NOR2X1 U15716 ( .A(conv_3[250]), .B(n28800), .Y(n29119) );
  NOR2X1 U15717 ( .A(conv_3[145]), .B(n33463), .Y(n33464) );
  NOR2X1 U15718 ( .A(conv_1[430]), .B(n29221), .Y(n29223) );
  NOR2X1 U15719 ( .A(conv_3[370]), .B(n33830), .Y(n33831) );
  NOR2X1 U15720 ( .A(conv_2[40]), .B(n33585), .Y(n33586) );
  NOR2X1 U15721 ( .A(n31252), .B(n31304), .Y(n31258) );
  NOR2X1 U15722 ( .A(conv_1[251]), .B(n26970), .Y(n26972) );
  NOR2X1 U15723 ( .A(n33636), .B(n35324), .Y(n27089) );
  NOR2X1 U15724 ( .A(conv_2[250]), .B(n33195), .Y(n33194) );
  NOR2X1 U15725 ( .A(conv_1[26]), .B(n30586), .Y(n30587) );
  NOR2X1 U15726 ( .A(n18203), .B(n18202), .Y(n25623) );
  NOR2X1 U15727 ( .A(n35135), .B(n24704), .Y(n18364) );
  NOR2X1 U15728 ( .A(ns[0]), .B(ns[1]), .Y(n20618) );
  NOR2X1 U15729 ( .A(n35162), .B(n35161), .Y(n35247) );
  NOR2X1 U15730 ( .A(n35201), .B(n26274), .Y(n26269) );
  AND4X2 U15731 ( .A(n21631), .B(n21630), .C(n21629), .D(n21628), .Y(n21632)
         );
  NOR2X1 U15732 ( .A(n20538), .B(n22713), .Y(n21382) );
  NOR2X1 U15733 ( .A(n20954), .B(n20953), .Y(n21028) );
  NOR2X1 U15734 ( .A(n35068), .B(n28575), .Y(n26206) );
  AND4X2 U15735 ( .A(n21590), .B(n21589), .C(n21588), .D(n21587), .Y(n21591)
         );
  NOR2X1 U15736 ( .A(n26023), .B(n26022), .Y(n26024) );
  NOR2X1 U15737 ( .A(n22716), .B(n28820), .Y(n22719) );
  NOR2X1 U15738 ( .A(n22550), .B(n30232), .Y(n20757) );
  NOR2X1 U15739 ( .A(n19401), .B(n33054), .Y(n19769) );
  AND4X2 U15740 ( .A(n21489), .B(n21488), .C(n21487), .D(n21486), .Y(n21490)
         );
  NOR2X1 U15741 ( .A(n16668), .B(n32256), .Y(n19526) );
  NOR2X1 U15742 ( .A(conv_3[24]), .B(n30199), .Y(n31252) );
  NOR2X1 U15743 ( .A(n31547), .B(n35823), .Y(n35829) );
  NOR2X1 U15744 ( .A(n31955), .B(n31967), .Y(n31974) );
  NOR2X1 U15745 ( .A(n30137), .B(n35884), .Y(n30148) );
  NOR2X1 U15746 ( .A(conv_1[70]), .B(n33635), .Y(n33636) );
  NOR2X1 U15747 ( .A(n27307), .B(n27311), .Y(n35295) );
  NOR2X1 U15748 ( .A(n35590), .B(n35593), .Y(n31227) );
  NOR2X1 U15749 ( .A(n29235), .B(n29240), .Y(n29215) );
  NOR2X1 U15750 ( .A(n33386), .B(n34775), .Y(n29298) );
  NOR2X1 U15751 ( .A(n35927), .B(n35930), .Y(n29928) );
  NOR2X1 U15752 ( .A(n33473), .B(n32130), .Y(n32128) );
  NOR2X1 U15753 ( .A(n35825), .B(n35821), .Y(n33960) );
  NOR2X1 U15754 ( .A(n22612), .B(n33134), .Y(n19773) );
  NOR2X1 U15755 ( .A(n22612), .B(n33985), .Y(n20761) );
  NOR2X1 U15756 ( .A(n28941), .B(n28936), .Y(n36066) );
  NOR2X1 U15757 ( .A(n31659), .B(n31655), .Y(n31649) );
  NOR2X1 U15758 ( .A(n32099), .B(n32095), .Y(n35672) );
  NOR2X1 U15759 ( .A(conv_2[219]), .B(n28667), .Y(n30430) );
  NOR2X1 U15760 ( .A(conv_2[474]), .B(n30901), .Y(n27881) );
  NOR2X1 U15761 ( .A(n31530), .B(n31529), .Y(n32059) );
  NOR2X1 U15762 ( .A(n36246), .B(n21388), .Y(n20542) );
  NOR2X1 U15763 ( .A(n28518), .B(n26285), .Y(n25355) );
  NOR2X1 U15764 ( .A(affine_2[41]), .B(n36225), .Y(n36227) );
  NOR2X1 U15765 ( .A(n25556), .B(n28479), .Y(n25012) );
  NOR2X1 U15766 ( .A(n26575), .B(n24708), .Y(n24713) );
  NOR2X1 U15767 ( .A(n35982), .B(n35983), .Y(n35981) );
  NOR2X1 U15768 ( .A(n27665), .B(n27670), .Y(n27672) );
  NOR2X1 U15769 ( .A(n21662), .B(n26039), .Y(n20303) );
  NOR2X1 U15770 ( .A(conv_3[339]), .B(n27590), .Y(n31955) );
  NOR2X1 U15771 ( .A(n34928), .B(n28467), .Y(n24701) );
  NOR2X1 U15772 ( .A(n26401), .B(n28349), .Y(n22675) );
  NOR2X1 U15773 ( .A(n25477), .B(n28349), .Y(n25486) );
  NOR2X1 U15774 ( .A(n31162), .B(n31166), .Y(n31179) );
  NOR2X1 U15775 ( .A(conv_2[54]), .B(n28713), .Y(n28712) );
  NOR2X1 U15776 ( .A(conv_3[204]), .B(n28838), .Y(n31849) );
  NOR2X1 U15777 ( .A(n35135), .B(n26549), .Y(n22699) );
  NOR2X1 U15778 ( .A(n36040), .B(n21536), .Y(n20843) );
  NOR2X1 U15779 ( .A(n21768), .B(n20320), .Y(n21760) );
  NOR2X1 U15780 ( .A(n29597), .B(n26085), .Y(n26031) );
  NOR2X1 U15781 ( .A(n26400), .B(n28577), .Y(n25389) );
  NOR2X1 U15782 ( .A(n28024), .B(n28023), .Y(n28767) );
  NOR2X1 U15783 ( .A(n22756), .B(n22755), .Y(n28554) );
  NOR2X1 U15784 ( .A(n21944), .B(n29425), .Y(n21812) );
  NOR2X1 U15785 ( .A(n33898), .B(n22008), .Y(n20552) );
  NOR2X1 U15786 ( .A(n19767), .B(n21435), .Y(n20565) );
  NOR2X1 U15787 ( .A(n25988), .B(n25987), .Y(n25991) );
  NOR2X1 U15788 ( .A(n33436), .B(n21953), .Y(n20060) );
  NOR2X1 U15789 ( .A(n21296), .B(n28277), .Y(n21298) );
  NOR2X1 U15790 ( .A(n36246), .B(n21357), .Y(n20481) );
  NOR2X1 U15791 ( .A(n22319), .B(n22318), .Y(n28643) );
  NOR2X1 U15792 ( .A(conv_3[489]), .B(n27616), .Y(n31547) );
  NOR2X1 U15793 ( .A(conv_2[114]), .B(n28682), .Y(n30137) );
  NOR2X1 U15794 ( .A(n21245), .B(n28479), .Y(n20505) );
  NOR2X1 U15795 ( .A(conv_2[414]), .B(n33689), .Y(n33690) );
  NOR2X1 U15796 ( .A(n33447), .B(n35591), .Y(n35589) );
  NOR2X1 U15797 ( .A(n32102), .B(n33478), .Y(n33007) );
  NOR2X1 U15798 ( .A(n33768), .B(n31121), .Y(n28667) );
  NOR2X1 U15799 ( .A(n23322), .B(n23326), .Y(n23316) );
  NOR2X1 U15800 ( .A(n27832), .B(n27831), .Y(n33619) );
  NOR2X1 U15801 ( .A(n36246), .B(n21313), .Y(n20476) );
  NOR2X1 U15802 ( .A(n18267), .B(n18266), .Y(n25576) );
  NOR2X1 U15803 ( .A(n22744), .B(n21688), .Y(n20320) );
  NOR2X1 U15804 ( .A(n19901), .B(n19900), .Y(n21662) );
  NOR2X1 U15805 ( .A(n19557), .B(n19556), .Y(n21433) );
  NOR2X1 U15806 ( .A(n29390), .B(n29394), .Y(n34291) );
  NOR2X1 U15807 ( .A(n35157), .B(n26473), .Y(n24844) );
  NOR2X1 U15808 ( .A(n22742), .B(n22741), .Y(n28579) );
  NOR2X1 U15809 ( .A(n18456), .B(n18455), .Y(n35041) );
  NOR2X1 U15810 ( .A(n22988), .B(n22992), .Y(n22993) );
  NOR2X1 U15811 ( .A(n35126), .B(n25123), .Y(n18612) );
  NOR2X1 U15812 ( .A(n36244), .B(n35133), .Y(n25701) );
  NOR2X1 U15813 ( .A(n28551), .B(n35070), .Y(n18560) );
  NOR2X1 U15814 ( .A(n19347), .B(n19346), .Y(n21290) );
  NOR2X1 U15815 ( .A(n20910), .B(n20909), .Y(n25963) );
  NOR2X1 U15816 ( .A(n22545), .B(n22544), .Y(n28442) );
  NOR2X1 U15817 ( .A(n19341), .B(n19340), .Y(n21285) );
  NOR2X1 U15818 ( .A(n27874), .B(n27873), .Y(n27886) );
  NOR2X1 U15819 ( .A(n25899), .B(n25892), .Y(n25896) );
  NOR2X1 U15820 ( .A(n21331), .B(n21329), .Y(n21343) );
  NOR2X1 U15821 ( .A(n21643), .B(n21639), .Y(n21642) );
  NOR2X1 U15822 ( .A(n22524), .B(n22523), .Y(n28519) );
  NOR2X1 U15823 ( .A(n29246), .B(n27259), .Y(n25260) );
  NOR2X1 U15824 ( .A(n18936), .B(n31016), .Y(n27910) );
  NOR2X1 U15825 ( .A(n16668), .B(n27362), .Y(n22769) );
  NOR2X1 U15826 ( .A(n31210), .B(n31215), .Y(n31205) );
  NOR2X1 U15827 ( .A(n25940), .B(n21863), .Y(n25943) );
  NOR2X1 U15828 ( .A(conv_2[8]), .B(n33568), .Y(n33569) );
  NOR2X1 U15829 ( .A(n29358), .B(n35471), .Y(n31280) );
  NOR2X1 U15830 ( .A(n27601), .B(n29823), .Y(n27172) );
  NOR2X1 U15831 ( .A(conv_1[24]), .B(n27609), .Y(n27608) );
  NOR2X1 U15832 ( .A(n31785), .B(n31790), .Y(n31798) );
  NOR2X1 U15833 ( .A(n22837), .B(n22842), .Y(n22832) );
  NOR2X1 U15834 ( .A(n34239), .B(n34243), .Y(n30077) );
  NOR2X1 U15835 ( .A(n26778), .B(n26777), .Y(n26790) );
  NOR2X1 U15836 ( .A(n31745), .B(n31749), .Y(n31751) );
  NOR2X1 U15837 ( .A(conv_3[457]), .B(n33776), .Y(n33777) );
  NOR2X1 U15838 ( .A(n29973), .B(n29972), .Y(n35527) );
  NOR2X1 U15839 ( .A(n31679), .B(n31684), .Y(n33743) );
  NOR2X1 U15840 ( .A(n26087), .B(n22014), .Y(n22020) );
  NOR2X1 U15841 ( .A(n36246), .B(n20553), .Y(n21418) );
  NOR2X1 U15842 ( .A(conv_3[322]), .B(n33839), .Y(n33840) );
  NOR2X1 U15843 ( .A(n33717), .B(n28959), .Y(n28958) );
  NOR2X1 U15844 ( .A(n35621), .B(n35625), .Y(n31413) );
  NOR2X1 U15845 ( .A(n18286), .B(n29086), .Y(n18288) );
  NOR2X1 U15846 ( .A(n32649), .B(n31597), .Y(n31596) );
  NOR2X1 U15847 ( .A(n18232), .B(n18231), .Y(n25522) );
  NOR2X1 U15848 ( .A(n18273), .B(n18272), .Y(n25575) );
  NOR2X1 U15849 ( .A(n18325), .B(n18324), .Y(n25556) );
  NOR2X1 U15850 ( .A(n21880), .B(n21358), .Y(n25899) );
  NOR2X1 U15851 ( .A(n21359), .B(n21358), .Y(n21360) );
  NOR2X1 U15852 ( .A(n19938), .B(n19937), .Y(n21560) );
  NOR2X1 U15853 ( .A(n18222), .B(n18221), .Y(n25587) );
  NOR2X1 U15854 ( .A(n21148), .B(n21358), .Y(n21149) );
  NOR2X1 U15855 ( .A(n24039), .B(n19918), .Y(n19920) );
  NOR2X1 U15856 ( .A(n24039), .B(n31130), .Y(n22592) );
  NOR2X1 U15857 ( .A(n21866), .B(n22713), .Y(n25940) );
  NOR2X1 U15858 ( .A(n18750), .B(n31858), .Y(n19304) );
  NOR2X1 U15859 ( .A(n18750), .B(n27325), .Y(n22570) );
  NOR2X1 U15860 ( .A(n18750), .B(n27321), .Y(n22554) );
  NOR2X1 U15861 ( .A(n18564), .B(n18563), .Y(n26223) );
  NOR2X1 U15862 ( .A(n18275), .B(n18274), .Y(n25583) );
  NOR2X1 U15863 ( .A(n18341), .B(n18340), .Y(n25604) );
  NOR2X1 U15864 ( .A(n22550), .B(n29668), .Y(n19363) );
  NOR2X1 U15865 ( .A(n18427), .B(n18426), .Y(n25205) );
  NOR2X1 U15866 ( .A(n36244), .B(n16755), .Y(n25795) );
  NOR2X1 U15867 ( .A(n22765), .B(n16661), .Y(n21833) );
  NOR2X1 U15868 ( .A(n35240), .B(n25123), .Y(n22245) );
  NOR2X1 U15869 ( .A(n18321), .B(n35381), .Y(n19922) );
  NOR2X1 U15870 ( .A(n19401), .B(n35722), .Y(n19403) );
  NOR2X1 U15871 ( .A(n19401), .B(n29485), .Y(n20854) );
  NOR2X1 U15872 ( .A(n19401), .B(n34160), .Y(n19574) );
  NOR2X1 U15873 ( .A(n19401), .B(n35277), .Y(n22486) );
  NOR2X1 U15874 ( .A(n22546), .B(n23450), .Y(n22614) );
  NOR2X1 U15875 ( .A(n22546), .B(n24924), .Y(n22548) );
  NOR2X1 U15876 ( .A(n18566), .B(n18565), .Y(n35085) );
  NOR2X1 U15877 ( .A(n34992), .B(n35231), .Y(n35184) );
  NOR2X1 U15878 ( .A(n27841), .B(n21953), .Y(n21958) );
  NOR2X1 U15879 ( .A(n22740), .B(n27099), .Y(n19895) );
  NOR2X1 U15880 ( .A(n36244), .B(n34982), .Y(n22244) );
  NOR2X1 U15881 ( .A(n35541), .B(n27220), .Y(n29973) );
  NOR2X1 U15882 ( .A(n35379), .B(n23439), .Y(n23444) );
  NOR2X1 U15883 ( .A(n33580), .B(n27771), .Y(n27775) );
  NOR2X1 U15884 ( .A(n35275), .B(n26505), .Y(n27334) );
  NOR2X1 U15885 ( .A(n35660), .B(n26526), .Y(n28831) );
  NOR2X1 U15886 ( .A(n35365), .B(n23593), .Y(n33193) );
  NOR2X1 U15887 ( .A(n16668), .B(n34311), .Y(n22731) );
  NOR2X1 U15888 ( .A(n22459), .B(n22458), .Y(n28502) );
  NOR2X1 U15889 ( .A(n18673), .B(n18672), .Y(n26280) );
  NOR2X1 U15890 ( .A(conv_1[397]), .B(n27639), .Y(n29358) );
  NOR2X1 U15891 ( .A(conv_1[292]), .B(n23170), .Y(n22826) );
  NOR2X1 U15892 ( .A(n36246), .B(n28479), .Y(n34903) );
  NOR2X1 U15893 ( .A(conv_1[367]), .B(n27576), .Y(n27575) );
  NOR2X1 U15894 ( .A(conv_3[157]), .B(n29749), .Y(n32248) );
  NOR2X1 U15895 ( .A(conv_3[502]), .B(n27629), .Y(n32065) );
  NOR2X1 U15896 ( .A(conv_2[68]), .B(n30118), .Y(n30120) );
  NOR2X1 U15897 ( .A(conv_1[201]), .B(n23680), .Y(n23681) );
  NOR2X1 U15898 ( .A(n33176), .B(n33088), .Y(n23134) );
  NOR2X1 U15899 ( .A(n31932), .B(n31931), .Y(n31939) );
  NOR2X1 U15900 ( .A(n30178), .B(n30183), .Y(n35869) );
  NOR2X1 U15901 ( .A(n36246), .B(n21172), .Y(n20433) );
  NOR2X1 U15902 ( .A(n22717), .B(n23398), .Y(n19897) );
  NOR2X1 U15903 ( .A(n22612), .B(n23155), .Y(n19915) );
  NOR2X1 U15904 ( .A(n28899), .B(n28903), .Y(n29947) );
  NOR2X1 U15905 ( .A(n36246), .B(n20513), .Y(n21331) );
  NOR2X1 U15906 ( .A(n36246), .B(n21879), .Y(n25892) );
  NOR2X1 U15907 ( .A(conv_2[381]), .B(n33415), .Y(n33416) );
  NOR2X1 U15908 ( .A(n31877), .B(n31881), .Y(n31890) );
  NOR2X1 U15909 ( .A(n34259), .B(n29383), .Y(n25274) );
  NOR2X1 U15910 ( .A(n32017), .B(n27764), .Y(n31180) );
  NOR2X1 U15911 ( .A(n26374), .B(n35241), .Y(n19179) );
  NOR2X1 U15912 ( .A(n29830), .B(n23296), .Y(n34626) );
  NOR2X1 U15913 ( .A(n35068), .B(n35198), .Y(n18556) );
  NOR2X1 U15914 ( .A(n24039), .B(n33693), .Y(n18265) );
  NOR2X1 U15915 ( .A(n24039), .B(n32015), .Y(n18583) );
  NOR2X1 U15916 ( .A(n24039), .B(n27808), .Y(n18238) );
  NOR2X1 U15917 ( .A(n18750), .B(n34393), .Y(n18477) );
  NOR2X1 U15918 ( .A(n18750), .B(n27029), .Y(n19840) );
  NOR2X1 U15919 ( .A(n18750), .B(n28679), .Y(n18242) );
  NOR2X1 U15920 ( .A(n22716), .B(n22571), .Y(n22573) );
  NOR2X1 U15921 ( .A(n21931), .B(n21688), .Y(n20810) );
  NOR2X1 U15922 ( .A(n22550), .B(n29908), .Y(n18339) );
  NOR2X1 U15923 ( .A(n22550), .B(n31442), .Y(n18581) );
  NOR2X1 U15924 ( .A(n34600), .B(n19044), .Y(n28137) );
  NOR2X1 U15925 ( .A(n18321), .B(n34362), .Y(n20896) );
  NOR2X1 U15926 ( .A(n18321), .B(n29188), .Y(n18323) );
  NOR2X1 U15927 ( .A(n32316), .B(n29747), .Y(n32284) );
  NOR2X1 U15928 ( .A(n18777), .B(n29902), .Y(n18230) );
  NOR2X1 U15929 ( .A(n18777), .B(n30066), .Y(n18308) );
  NOR2X1 U15930 ( .A(n19274), .B(n19273), .Y(n21243) );
  NOR2X1 U15931 ( .A(n35463), .B(n19153), .Y(n33181) );
  NOR2X1 U15932 ( .A(n22740), .B(n34221), .Y(n18411) );
  NOR2X1 U15933 ( .A(n22740), .B(n31237), .Y(n18515) );
  NOR2X1 U15934 ( .A(n35441), .B(n24319), .Y(n26364) );
  NOR2X1 U15935 ( .A(n34132), .B(n27741), .Y(n27747) );
  NOR2X1 U15936 ( .A(n34211), .B(n28133), .Y(n28892) );
  NOR2X1 U15937 ( .A(n35404), .B(n22299), .Y(n33187) );
  NOR2X1 U15938 ( .A(n33787), .B(n35775), .Y(n35767) );
  NOR2X1 U15939 ( .A(conv_3[96]), .B(n33741), .Y(n33742) );
  NOR2X1 U15940 ( .A(n33593), .B(n35862), .Y(n27728) );
  NOR2X1 U15941 ( .A(conv_3[321]), .B(n28759), .Y(n31907) );
  NOR2X1 U15942 ( .A(n28696), .B(n19173), .Y(n30202) );
  NOR2X1 U15943 ( .A(n22612), .B(n22816), .Y(n19936) );
  NOR2X1 U15944 ( .A(n22717), .B(n30075), .Y(n18220) );
  NOR2X1 U15945 ( .A(n22612), .B(n30159), .Y(n18306) );
  NOR2X1 U15946 ( .A(n34125), .B(n34128), .Y(n33805) );
  NOR2X1 U15947 ( .A(n25247), .B(n22269), .Y(n34259) );
  NOR2X1 U15948 ( .A(affine_2[21]), .B(n36215), .Y(n36217) );
  NOR2X1 U15949 ( .A(n28290), .B(n20755), .Y(n21736) );
  NOR2X1 U15950 ( .A(n32017), .B(n31418), .Y(n35599) );
  NOR2X1 U15951 ( .A(n29830), .B(n22269), .Y(n35982) );
  NOR2X1 U15952 ( .A(n19221), .B(n19181), .Y(n25399) );
  AOI222XL U15953 ( .A0(conv_3[5]), .A1(n34379), .B0(n32996), .B1(n24370), 
        .C0(n28689), .C1(n28687), .Y(n31427) );
  NOR2X1 U15954 ( .A(n32017), .B(n27860), .Y(n35810) );
  NOR2X1 U15955 ( .A(n25247), .B(n33422), .Y(n27131) );
  NOR2X1 U15956 ( .A(n36244), .B(n24971), .Y(n25116) );
  NOR2X1 U15957 ( .A(n22550), .B(n32289), .Y(n19282) );
  NOR2X1 U15958 ( .A(n22550), .B(n23227), .Y(n18503) );
  NOR2X1 U15959 ( .A(n33096), .B(n29139), .Y(n29512) );
  NOR2X1 U15960 ( .A(n22765), .B(n28277), .Y(n21464) );
  NOR2X1 U15961 ( .A(n18776), .B(n22150), .Y(n18492) );
  NOR2X1 U15962 ( .A(n32887), .B(n18855), .Y(n33166) );
  NOR2X1 U15963 ( .A(conv_3[455]), .B(n35795), .Y(n35798) );
  NOR2X1 U15964 ( .A(conv_3[426]), .B(n33786), .Y(n33787) );
  NOR2X1 U15965 ( .A(n32025), .B(n32024), .Y(n32031) );
  NOR2X1 U15966 ( .A(conv_2[35]), .B(n33592), .Y(n33593) );
  NOR2X1 U15967 ( .A(conv_2[516]), .B(n33577), .Y(n33578) );
  NOR2X1 U15968 ( .A(conv_1[230]), .B(n33183), .Y(n33182) );
  NOR2X1 U15969 ( .A(conv_1[185]), .B(n33189), .Y(n33188) );
  NOR2X1 U15970 ( .A(conv_2[276]), .B(n18956), .Y(n28024) );
  NOR2X1 U15971 ( .A(n35750), .B(n31967), .Y(n35753) );
  NOR2X1 U15972 ( .A(conv_3[35]), .B(n35582), .Y(n35585) );
  ADDFX2 U15973 ( .A(conv_3[126]), .B(n35622), .CI(n32662), .CO(n35623), .S(
        n32663) );
  NOR2X1 U15974 ( .A(n22612), .B(n22881), .Y(n18497) );
  NOR2X1 U15975 ( .A(n36246), .B(n21242), .Y(n19280) );
  NOR2X1 U15976 ( .A(n32017), .B(n19108), .Y(n35732) );
  NOR2X1 U15977 ( .A(n27538), .B(n22262), .Y(n35344) );
  NOR2X1 U15978 ( .A(n28602), .B(n23290), .Y(n23341) );
  NOR2X1 U15979 ( .A(n29830), .B(n27532), .Y(n34529) );
  NOR2X1 U15980 ( .A(n25247), .B(n27532), .Y(n35463) );
  NOR2X1 U15981 ( .A(n23426), .B(n23425), .Y(n30695) );
  NOR2X1 U15982 ( .A(n22546), .B(n31718), .Y(n18554) );
  NOR2X1 U15983 ( .A(n25247), .B(n23296), .Y(n34044) );
  NOR2X1 U15984 ( .A(n29455), .B(n28149), .Y(n28258) );
  NOR2X1 U15985 ( .A(n33979), .B(n19114), .Y(n30858) );
  NOR2X1 U15986 ( .A(conv_2[500]), .B(n31017), .Y(n18936) );
  NOR2X1 U15987 ( .A(conv_3[335]), .B(n35746), .Y(n35750) );
  NOR2X1 U15988 ( .A(conv_1[470]), .B(n33162), .Y(n33161) );
  NOR2X1 U15989 ( .A(conv_2[410]), .B(n33377), .Y(n33380) );
  NOR2X1 U15990 ( .A(conv_1[259]), .B(n33215), .Y(n33214) );
  NOR2X1 U15991 ( .A(n29830), .B(n22257), .Y(n29831) );
  NOR2X1 U15992 ( .A(n27644), .B(n35858), .Y(n27642) );
  NOR2X1 U15993 ( .A(n24318), .B(n24317), .Y(n30283) );
  NOR2X1 U15994 ( .A(n26513), .B(n26512), .Y(n26922) );
  NOR2X1 U15995 ( .A(n31691), .B(n27860), .Y(n19020) );
  NOR2X1 U15996 ( .A(n22164), .B(n22163), .Y(n26152) );
  NOR2X1 U15997 ( .A(n32959), .B(n17143), .Y(n16773) );
  NOR2X1 U15998 ( .A(n35500), .B(n27898), .Y(n23642) );
  NOR2X1 U15999 ( .A(n17013), .B(n17012), .Y(n17015) );
  NOR2X1 U16000 ( .A(conv_1[515]), .B(n27261), .Y(n24913) );
  NOR2X1 U16001 ( .A(n35856), .B(n22269), .Y(n24296) );
  NOR2X1 U16002 ( .A(n25247), .B(n22257), .Y(n23923) );
  NOR2X1 U16003 ( .A(n17969), .B(n28611), .Y(DP_OP_5171J1_127_4278_n89) );
  NOR2X1 U16004 ( .A(n17969), .B(n28398), .Y(DP_OP_5170J1_126_4278_n89) );
  NOR2X1 U16005 ( .A(n19652), .B(n28211), .Y(DP_OP_5169J1_125_4278_n89) );
  NOR2X1 U16006 ( .A(n33403), .B(n34715), .Y(n24346) );
  NOR2X1 U16007 ( .A(n33403), .B(n34522), .Y(n22980) );
  NOR2X1 U16008 ( .A(n33403), .B(n23296), .Y(n24428) );
  NOR2X1 U16009 ( .A(n28664), .B(n28663), .Y(n28877) );
  NOR2X1 U16010 ( .A(n27687), .B(n27686), .Y(n28853) );
  NOR2X1 U16011 ( .A(n34164), .B(n31455), .Y(n31454) );
  NOR2X1 U16012 ( .A(n35858), .B(n27532), .Y(n23078) );
  NOR2X1 U16013 ( .A(n35856), .B(n32016), .Y(n24449) );
  NOR2X1 U16014 ( .A(n32017), .B(n22257), .Y(n35639) );
  NOR2X1 U16015 ( .A(n35500), .B(n27848), .Y(n23438) );
  NOR2X1 U16016 ( .A(n27644), .B(n31691), .Y(n24260) );
  NOR2X1 U16017 ( .A(n32017), .B(n28948), .Y(n35622) );
  NOR2X1 U16018 ( .A(n22877), .B(n22876), .Y(n31666) );
  NOR2X1 U16019 ( .A(n23591), .B(n23590), .Y(n23976) );
  NOR2X1 U16020 ( .A(n31691), .B(n24021), .Y(n24026) );
  NOR2X1 U16021 ( .A(n16835), .B(n16834), .Y(n16836) );
  NOR2X1 U16022 ( .A(n30242), .B(n18971), .Y(n30112) );
  NOR2X1 U16023 ( .A(n35498), .B(n22257), .Y(n22434) );
  NOR2X1 U16024 ( .A(n35498), .B(n24021), .Y(n24272) );
  NOR2X1 U16025 ( .A(n29426), .B(n33020), .Y(n23730) );
  NOR2X1 U16026 ( .A(n17144), .B(n19182), .Y(n17068) );
  NOR2X1 U16027 ( .A(n23550), .B(n23549), .Y(n24364) );
  NOR2X1 U16028 ( .A(n35856), .B(n23504), .Y(n23234) );
  NOR2X1 U16029 ( .A(n32017), .B(n27532), .Y(n34164) );
  NOR2X1 U16030 ( .A(n33988), .B(n35858), .Y(n27706) );
  NOR2X1 U16031 ( .A(n35856), .B(n23296), .Y(n23112) );
  NOR2X1 U16032 ( .A(n27848), .B(n32017), .Y(n35653) );
  NOR2X1 U16033 ( .A(n23768), .B(n23767), .Y(n26945) );
  NOR2X1 U16034 ( .A(n32729), .B(n17143), .Y(n16826) );
  NOR2X1 U16035 ( .A(n35856), .B(n33429), .Y(n27685) );
  NOR2X1 U16036 ( .A(n35498), .B(n28948), .Y(n23646) );
  NOR2X1 U16037 ( .A(n18997), .B(n27860), .Y(n30780) );
  NOR2X1 U16038 ( .A(n35856), .B(n28660), .Y(n28662) );
  NOR2X1 U16039 ( .A(n19643), .B(n19652), .Y(n19646) );
  NOR2X1 U16040 ( .A(n19622), .B(n19652), .Y(n19625) );
  NOR2X1 U16041 ( .A(n35500), .B(n33429), .Y(n22218) );
  NOR2X1 U16042 ( .A(n18997), .B(n34715), .Y(n30794) );
  NOR2X1 U16043 ( .A(n35498), .B(n27532), .Y(n23194) );
  NOR2X1 U16044 ( .A(n19182), .B(n17391), .Y(n17454) );
  NOR2X1 U16045 ( .A(n35498), .B(n34426), .Y(n26749) );
  NOR2X1 U16046 ( .A(n35498), .B(n27799), .Y(n27327) );
  NOR2X1 U16047 ( .A(n29426), .B(n19108), .Y(n23486) );
  NOR2X1 U16048 ( .A(n35500), .B(n27764), .Y(n27386) );
  NOR2X1 U16049 ( .A(n33403), .B(n27898), .Y(n30581) );
  NOR2X1 U16050 ( .A(n33403), .B(n19215), .Y(n24514) );
  NOR2X1 U16051 ( .A(n27848), .B(n35853), .Y(n27416) );
  NOR2X1 U16052 ( .A(n35498), .B(n33422), .Y(n23423) );
  NOR2X1 U16053 ( .A(n31691), .B(n28948), .Y(n23690) );
  NOR2X1 U16054 ( .A(n34714), .B(n22931), .Y(n22932) );
  NOR2X1 U16055 ( .A(n27624), .B(n27623), .Y(n29631) );
  NOR2X1 U16056 ( .A(n22181), .B(n22180), .Y(n29959) );
  AOI222XL U16057 ( .A0(n30401), .A1(conv_2[377]), .B0(n30401), .B1(n30400), 
        .C0(conv_2[377]), .C1(n30400), .Y(n23075) );
  AOI222XL U16058 ( .A0(n27289), .A1(conv_2[78]), .B0(n27289), .B1(n27288), 
        .C0(conv_2[78]), .C1(n27288), .Y(n23479) );
  NOR2X1 U16059 ( .A(n29429), .B(n29428), .Y(n30549) );
  NOR2X1 U16060 ( .A(n33403), .B(n27848), .Y(n24142) );
  NOR2X1 U16061 ( .A(n18997), .B(n23504), .Y(n23562) );
  NOR2X1 U16062 ( .A(n35498), .B(n27764), .Y(n30456) );
  NOR2X1 U16063 ( .A(n20601), .B(n17026), .Y(n17038) );
  NOR2X1 U16064 ( .A(n19652), .B(n19691), .Y(n19676) );
  NOR2X1 U16065 ( .A(n18997), .B(n24021), .Y(n24023) );
  NOR2X1 U16066 ( .A(n35856), .B(n22257), .Y(n29002) );
  NOR2X1 U16067 ( .A(n19192), .B(n19191), .Y(n24203) );
  NOR2X1 U16068 ( .A(n35853), .B(n24021), .Y(n30273) );
  NOR2X1 U16069 ( .A(n30536), .B(n29427), .Y(n29429) );
  NOR2X1 U16070 ( .A(n17969), .B(n19630), .Y(n19673) );
  NOR2X1 U16071 ( .A(n33403), .B(n27644), .Y(n27380) );
  NOR2X1 U16072 ( .A(n21536), .B(n19182), .Y(n17842) );
  NOR2X1 U16073 ( .A(n35856), .B(n31871), .Y(n28087) );
  NOR2X1 U16074 ( .A(n18913), .B(n23101), .Y(n23102) );
  NOR2X1 U16075 ( .A(n35498), .B(n33988), .Y(n26977) );
  NOR2X1 U16076 ( .A(n35498), .B(n27735), .Y(n27225) );
  NOR2X1 U16077 ( .A(n35498), .B(n29136), .Y(n23364) );
  NOR2X1 U16078 ( .A(n35856), .B(n33020), .Y(n27289) );
  NOR2X1 U16079 ( .A(n18997), .B(n29136), .Y(n30846) );
  NOR2X1 U16080 ( .A(n35564), .B(n35563), .Y(n35562) );
  NOR2X1 U16081 ( .A(n20726), .B(n17172), .Y(n17755) );
  NOR2X1 U16082 ( .A(n33403), .B(n19128), .Y(n26915) );
  NOR2X1 U16083 ( .A(n33403), .B(n26128), .Y(n27438) );
  NOR2X1 U16084 ( .A(n34703), .B(n29426), .Y(n29732) );
  NOR2X1 U16085 ( .A(n33403), .B(n33402), .Y(n33539) );
  NOR2X1 U16086 ( .A(n24490), .B(n24488), .Y(n24486) );
  NOR2X1 U16087 ( .A(n19416), .B(n16707), .Y(n17753) );
  NOR2X1 U16088 ( .A(n19214), .B(n24525), .Y(n19215) );
  NOR2X1 U16089 ( .A(n27900), .B(n27899), .Y(n30394) );
  NOR2X1 U16090 ( .A(n18913), .B(n24445), .Y(n30306) );
  NOR2X1 U16091 ( .A(n28073), .B(n28072), .Y(n29420) );
  NOR2X1 U16092 ( .A(n22269), .B(n22270), .Y(n33860) );
  NOR2X1 U16093 ( .A(n18997), .B(n28721), .Y(n30575) );
  NOR2X1 U16094 ( .A(n34703), .B(n35853), .Y(n27082) );
  NOR2X1 U16095 ( .A(n33403), .B(n27532), .Y(n19149) );
  NOR2X1 U16096 ( .A(n18997), .B(n32016), .Y(n30852) );
  NOR2X1 U16097 ( .A(n35498), .B(n27860), .Y(n26952) );
  NOR2X1 U16098 ( .A(n26509), .B(n18997), .Y(n30824) );
  NOR2X1 U16099 ( .A(n29426), .B(n27799), .Y(n29720) );
  NOR2X1 U16100 ( .A(n33403), .B(n34703), .Y(n23970) );
  NOR2X1 U16101 ( .A(n35856), .B(n27764), .Y(n29644) );
  NOR2X1 U16102 ( .A(n29426), .B(n27532), .Y(n19192) );
  NOR2X1 U16103 ( .A(n18997), .B(n23296), .Y(n30818) );
  NOR2X1 U16104 ( .A(n33403), .B(n27215), .Y(n27373) );
  NOR2X1 U16105 ( .A(n30536), .B(n31108), .Y(n30525) );
  NOR2X1 U16106 ( .A(n33403), .B(n23463), .Y(n23466) );
  NOR2X1 U16107 ( .A(n29426), .B(n28948), .Y(n35570) );
  NOR2X1 U16108 ( .A(n27764), .B(n23256), .Y(n27062) );
  NOR2X1 U16109 ( .A(n24672), .B(n24670), .Y(n24668) );
  NOR2X1 U16110 ( .A(n24559), .B(n24557), .Y(n24555) );
  NOR2X1 U16111 ( .A(n22897), .B(n34425), .Y(n22899) );
  NOR2X1 U16112 ( .A(n33401), .B(n33400), .Y(n33402) );
  NOR2X1 U16113 ( .A(n30536), .B(n31329), .Y(n30562) );
  NOR2X1 U16114 ( .A(n22916), .B(n33019), .Y(n22918) );
  NOR2X1 U16115 ( .A(n34522), .B(n23082), .Y(n34485) );
  NOR2X1 U16116 ( .A(n24277), .B(n24520), .Y(n29761) );
  OAI211X4 U16117 ( .A0(n20389), .A1(n18119), .B0(n18105), .C0(n18104), .Y(
        n18106) );
  NOR2X1 U16118 ( .A(n33403), .B(n28070), .Y(n30736) );
  NOR2X1 U16119 ( .A(n20755), .B(n18043), .Y(n17813) );
  NOR2X1 U16120 ( .A(n35853), .B(n31418), .Y(n24251) );
  NOR2X1 U16121 ( .A(n26207), .B(n18043), .Y(n17826) );
  NOR2X1 U16122 ( .A(n27848), .B(n18997), .Y(n30800) );
  NOR2X1 U16123 ( .A(n18286), .B(n35239), .Y(n17886) );
  NOR2X1 U16124 ( .A(n35853), .B(n27764), .Y(n27766) );
  NOR2X1 U16125 ( .A(n18286), .B(n28553), .Y(n17810) );
  NOR2X1 U16126 ( .A(n18286), .B(n28479), .Y(n17874) );
  NOR2X1 U16127 ( .A(n18997), .B(n35499), .Y(n30806) );
  NOR2X1 U16128 ( .A(n22740), .B(n34981), .Y(n17893) );
  NOR2X1 U16129 ( .A(n35856), .B(n19108), .Y(n24185) );
  NOR2X1 U16130 ( .A(n29426), .B(n22257), .Y(n29069) );
  NOR2X1 U16131 ( .A(n26509), .B(n35856), .Y(n23032) );
  NOR2X1 U16132 ( .A(n35159), .B(n22018), .Y(n17815) );
  NOR2X1 U16133 ( .A(n19902), .B(n26279), .Y(n17863) );
  NOR2X1 U16134 ( .A(n22716), .B(n34981), .Y(n17873) );
  NOR2X1 U16135 ( .A(n22717), .B(n28479), .Y(n17867) );
  NOR2X1 U16136 ( .A(n35853), .B(n28070), .Y(n29966) );
  NOR2X1 U16137 ( .A(n35159), .B(n19182), .Y(n17166) );
  NOR2X1 U16138 ( .A(n19247), .B(n19246), .Y(n20363) );
  NOR2X1 U16139 ( .A(n22716), .B(n26621), .Y(n17825) );
  NOR2X1 U16140 ( .A(n18997), .B(n34522), .Y(n30623) );
  NOR2X1 U16141 ( .A(n18997), .B(n27898), .Y(n30812) );
  NOR2X1 U16142 ( .A(n16715), .B(n26621), .Y(n17827) );
  NOR2X1 U16143 ( .A(n18925), .B(n18924), .Y(n30319) );
  NOR2X1 U16144 ( .A(n18997), .B(n23686), .Y(n30741) );
  NOR2X1 U16145 ( .A(n24524), .B(n24522), .Y(n24520) );
  NOR2X1 U16146 ( .A(n27620), .B(n31871), .Y(n30619) );
  NOR2X1 U16147 ( .A(n18913), .B(n27897), .Y(n30312) );
  NOR2X1 U16148 ( .A(n30536), .B(n30602), .Y(n33547) );
  NOR2X1 U16149 ( .A(n35272), .B(n34764), .Y(n24277) );
  NOR2X1 U16150 ( .A(n25074), .B(n25073), .Y(n25075) );
  NOR2X1 U16151 ( .A(n22429), .B(n23884), .Y(n30466) );
  OAI211X4 U16152 ( .A0(n20405), .A1(n18119), .B0(n18083), .C0(n18082), .Y(
        n18084) );
  NOR2X1 U16153 ( .A(n18913), .B(n34416), .Y(n23097) );
  NOR2X1 U16154 ( .A(n34703), .B(n23568), .Y(n34510) );
  NOR2X1 U16155 ( .A(n27799), .B(n23024), .Y(n34506) );
  NOR2X1 U16156 ( .A(conv_3[167]), .B(n35554), .Y(n35558) );
  NOR2X1 U16157 ( .A(n27644), .B(n19058), .Y(n28718) );
  NOR2X1 U16158 ( .A(n30536), .B(n30610), .Y(n30556) );
  NOR2X1 U16159 ( .A(n30536), .B(n31380), .Y(n30729) );
  NOR2X1 U16160 ( .A(n23792), .B(n24266), .Y(n23793) );
  NOR2X1 U16161 ( .A(n23943), .B(n23945), .Y(n23941) );
  NOR2X1 U16162 ( .A(n33429), .B(n24306), .Y(n34497) );
  NOR2X1 U16163 ( .A(n30536), .B(n35499), .Y(n29679) );
  NOR2X1 U16164 ( .A(n27620), .B(n25456), .Y(n25454) );
  NOR2X1 U16165 ( .A(n33423), .B(n32016), .Y(n30649) );
  NOR2X1 U16166 ( .A(n33989), .B(n34715), .Y(n22855) );
  NOR2X1 U16167 ( .A(n33423), .B(n35857), .Y(n26957) );
  NOR2X1 U16168 ( .A(n18913), .B(n22882), .Y(n34233) );
  NOR2X1 U16169 ( .A(n33989), .B(n24021), .Y(n23146) );
  NOR2X1 U16170 ( .A(n30536), .B(n27042), .Y(n30568) );
  NOR2X1 U16171 ( .A(n27898), .B(n33989), .Y(n22893) );
  NOR2X1 U16172 ( .A(n23831), .B(n18913), .Y(n35844) );
  NOR2X1 U16173 ( .A(n27531), .B(n19188), .Y(n19189) );
  NOR2X1 U16174 ( .A(n27848), .B(n33989), .Y(n34115) );
  NOR2X1 U16175 ( .A(n35272), .B(n33528), .Y(n27214) );
  NOR2X1 U16176 ( .A(n35272), .B(n33864), .Y(n19214) );
  NOR2X1 U16177 ( .A(n33423), .B(n33994), .Y(n30653) );
  NOR2X1 U16178 ( .A(n24940), .B(n24942), .Y(n27213) );
  INVX2 U16179 ( .A(n34476), .Y(n28660) );
  NOR2X1 U16180 ( .A(n35272), .B(n33428), .Y(n22215) );
  NOR2X1 U16181 ( .A(n30536), .B(n30837), .Y(n27513) );
  NOR2X1 U16182 ( .A(n33423), .B(n26509), .Y(n26695) );
  NOR2X1 U16183 ( .A(n27620), .B(n22269), .Y(n30611) );
  AOI211X2 U16184 ( .A0(n34827), .A1(n23090), .B0(n22214), .C0(n22213), .Y(
        n33429) );
  NOR2X1 U16185 ( .A(n33989), .B(n28070), .Y(n24209) );
  NOR2X1 U16186 ( .A(n33989), .B(n31418), .Y(n23832) );
  INVX2 U16187 ( .A(n34502), .Y(n23504) );
  NOR2X1 U16188 ( .A(n18913), .B(n33020), .Y(n23473) );
  NOR2X1 U16189 ( .A(n33422), .B(n33989), .Y(n22883) );
  NOR2X1 U16190 ( .A(n27483), .B(n27479), .Y(n23748) );
  NOR2X1 U16191 ( .A(n35857), .B(n27620), .Y(n31027) );
  INVX2 U16192 ( .A(n27691), .Y(n35857) );
  INVX2 U16193 ( .A(n34706), .Y(n34703) );
  NOR2X1 U16194 ( .A(n27620), .B(n28948), .Y(n30838) );
  NAND2X1 U16195 ( .A(n16725), .B(n28290), .Y(n18118) );
  BUFX2 U16196 ( .A(n22426), .Y(n28948) );
  NOR2X1 U16197 ( .A(n33989), .B(n34439), .Y(n34436) );
  INVX2 U16198 ( .A(n34422), .Y(n28721) );
  AOI21X2 U16199 ( .A0(n26470), .A1(n23089), .B0(n22256), .Y(n22257) );
  NOR2X1 U16200 ( .A(n36244), .B(n26479), .Y(n34921) );
  NOR2X1 U16201 ( .A(n36244), .B(n35241), .Y(n25766) );
  INVX2 U16202 ( .A(n34450), .Y(n26509) );
  NOR2X1 U16203 ( .A(n36244), .B(n35159), .Y(n23785) );
  NOR2X1 U16204 ( .A(n21095), .B(n28277), .Y(n21097) );
  INVX2 U16205 ( .A(n18172), .Y(n19008) );
  NOR2X1 U16206 ( .A(n19221), .B(n16721), .Y(n23276) );
  INVX2 U16207 ( .A(n19227), .Y(n19009) );
  INVX2 U16208 ( .A(n19416), .Y(n22021) );
  NOR2X1 U16209 ( .A(n26374), .B(n23052), .Y(n18475) );
  NOR2X1 U16210 ( .A(n36248), .B(counter[1]), .Y(n17988) );
  NOR2X1 U16211 ( .A(N18471), .B(n16721), .Y(n26172) );
  BUFX2 U16212 ( .A(n16722), .Y(n28290) );
  NOR2X1 U16213 ( .A(n28292), .B(n16715), .Y(n16709) );
  NOR2X1 U16214 ( .A(n19181), .B(n35159), .Y(n16746) );
  INVX2 U16215 ( .A(n22370), .Y(n19181) );
  BUFX8 U16216 ( .A(cursor[5]), .Y(n36244) );
  INVX4 U16217 ( .A(N18014), .Y(n19221) );
  NOR2XL U16218 ( .A(n18174), .B(n34891), .Y(n16967) );
  NOR2XL U16219 ( .A(n16669), .B(n16707), .Y(n17848) );
  NOR2XL U16220 ( .A(n22716), .B(n28814), .Y(n22622) );
  NOR2XL U16221 ( .A(n16715), .B(n33110), .Y(n19555) );
  NOR2XL U16222 ( .A(n17173), .B(n17172), .Y(n17847) );
  NOR2XL U16223 ( .A(n17165), .B(n17172), .Y(n17854) );
  NOR2XL U16224 ( .A(n22716), .B(n34561), .Y(n22492) );
  NOR2XL U16225 ( .A(n16715), .B(n35284), .Y(n22462) );
  NOR2XL U16226 ( .A(n16715), .B(n23375), .Y(n22711) );
  NOR2XL U16227 ( .A(n22716), .B(n32226), .Y(n18657) );
  BUFX2 U16228 ( .A(n16735), .Y(n18127) );
  OAI221X1 U16229 ( .A0(n18133), .A1(n24571), .B0(n18132), .B1(n18128), .C0(
        n28611), .Y(n28610) );
  AOI222XL U16230 ( .A0(n28087), .A1(conv_2[288]), .B0(n28087), .B1(n28086), 
        .C0(conv_2[288]), .C1(n28086), .Y(n28088) );
  NOR2X1 U16231 ( .A(counter[2]), .B(n16675), .Y(n19005) );
  ADDFXL U16232 ( .A(n17921), .B(affine_1[7]), .CI(n17920), .CO(
        DP_OP_5168J1_124_9881_n18), .S(DP_OP_5168J1_124_9881_n19) );
  XOR2XL U16233 ( .A(n33070), .B(DP_OP_5168J1_124_9881_n13), .Y(n33072) );
  ADDFXL U16234 ( .A(n17159), .B(n17158), .CI(n17157), .CO(
        DP_OP_5166J1_122_9881_n37), .S(DP_OP_5166J1_122_9881_n38) );
  NOR2XL U16235 ( .A(n29426), .B(n28721), .Y(n22113) );
  NOR2XL U16236 ( .A(n35858), .B(n22257), .Y(n29004) );
  AOI222XL U16237 ( .A0(n35009), .A1(n35008), .B0(n35009), .B1(n28303), .C0(
        n35008), .C1(n28303), .Y(n28362) );
  NOR2XL U16238 ( .A(n23696), .B(conv_1[530]), .Y(n22222) );
  NOR2XL U16239 ( .A(n29136), .B(n35500), .Y(n22298) );
  INVXL U16240 ( .A(n18321), .Y(n18240) );
  INVX2 U16241 ( .A(n27429), .Y(n35272) );
  INVX2 U16242 ( .A(n18782), .Y(n16670) );
  NOR2XL U16243 ( .A(n35498), .B(n35857), .Y(intadd_2_B_1_) );
  NAND2X1 U16244 ( .A(n36245), .B(N17708), .Y(n21830) );
  INVXL U16245 ( .A(n27990), .Y(n32016) );
  NAND2X2 U16246 ( .A(n28407), .B(n34827), .Y(n35239) );
  ADDFX2 U16247 ( .A(DP_OP_5167J1_123_9881_n21), .B(DP_OP_5167J1_123_9881_n17), 
        .CI(n25242), .CO(n33555), .S(n22197) );
  ADDFX2 U16248 ( .A(DP_OP_5166J1_122_9881_n43), .B(n20695), .CI(n20694), .CO(
        n20703), .S(n20696) );
  ADDFXL U16249 ( .A(conv_2[48]), .B(n27801), .CI(n27800), .CO(n29740), .S(
        n23029) );
  INVX4 U16250 ( .A(n16745), .Y(n28479) );
  NOR2XL U16251 ( .A(n31419), .B(n31420), .Y(n23902) );
  ADDFXL U16252 ( .A(conv_1[417]), .B(n35493), .CI(n34671), .CO(n34776), .S(
        n32688) );
  NOR2XL U16253 ( .A(n25247), .B(n28070), .Y(n35493) );
  ADDFXL U16254 ( .A(conv_1[325]), .B(n34259), .CI(n22926), .CO(n34258), .S(
        n22275) );
  ADDFXL U16255 ( .A(conv_1[248]), .B(n33663), .CI(n23835), .CO(n35411), .S(
        n23660) );
  ADDFXL U16256 ( .A(conv_1[157]), .B(n34044), .CI(n24312), .CO(n34043), .S(
        n24313) );
  ADDFXL U16257 ( .A(conv_1[130]), .B(n34292), .CI(n25447), .CO(n30450), .S(
        n23651) );
  ADDFXL U16258 ( .A(conv_1[9]), .B(n27278), .CI(n24537), .CO(n27279), .S(
        n22381) );
  ADDFXL U16259 ( .A(conv_2[156]), .B(n34626), .CI(n24530), .CO(n29863), .S(
        n23116) );
  ADDFXL U16260 ( .A(conv_2[128]), .B(n34344), .CI(n24361), .CO(n34343), .S(
        n24355) );
  NOR2XL U16261 ( .A(n32017), .B(n28070), .Y(n32557) );
  NOR2XL U16262 ( .A(n31615), .B(n31614), .Y(n31617) );
  NOR2XL U16263 ( .A(n31431), .B(n31430), .Y(n31433) );
  NOR2XL U16264 ( .A(n19221), .B(n35262), .Y(n19226) );
  NOR2XL U16265 ( .A(n23052), .B(n35262), .Y(n35258) );
  INVXL U16266 ( .A(n35641), .Y(n35630) );
  INVXL U16267 ( .A(n16734), .Y(n21944) );
  NOR2X2 U16268 ( .A(n36245), .B(n18286), .Y(n16734) );
  INVXL U16269 ( .A(n21954), .Y(n16669) );
  INVX2 U16270 ( .A(n22368), .Y(n18239) );
  INVX2 U16271 ( .A(n20978), .Y(n19902) );
  INVXL U16272 ( .A(n36042), .Y(n32656) );
  INVX2 U16273 ( .A(n36001), .Y(n16656) );
  OAI211XL U16274 ( .A0(n34789), .A1(n33911), .B0(n33468), .C0(n33910), .Y(
        n15564) );
  OAI2BB1XL U16275 ( .A0N(conv_1[235]), .A1N(n31128), .B0(n34276), .Y(n34275)
         );
  NOR2X1 U16276 ( .A(n35404), .B(n35405), .Y(n35403) );
  AOI21XL U16277 ( .A0(n26341), .A1(n26346), .B0(n26342), .Y(n32886) );
  NOR2BXL U16278 ( .AN(n35977), .B(n35978), .Y(n33978) );
  NOR2X1 U16279 ( .A(conv_3[386]), .B(n32197), .Y(n32199) );
  AOI32XL U16280 ( .A0(n35626), .A1(n28955), .A2(n28954), .B0(n31436), .B1(
        n28955), .Y(n15659) );
  NOR2X1 U16281 ( .A(n30586), .B(n33202), .Y(n27336) );
  NOR2X1 U16282 ( .A(n28172), .B(n36042), .Y(n28173) );
  NOR2BXL U16283 ( .AN(n35714), .B(n35715), .Y(n33226) );
  NOR2X1 U16284 ( .A(n32131), .B(n32130), .Y(n33724) );
  NOR2BXL U16285 ( .AN(n35964), .B(n35965), .Y(n32976) );
  AOI32XL U16286 ( .A0(n31013), .A1(n28710), .A2(n28709), .B0(n28708), .B1(
        n28710), .Y(n14859) );
  NAND2XL U16287 ( .A(n35891), .B(n30138), .Y(n34364) );
  NOR2X1 U16288 ( .A(n33812), .B(n30924), .Y(n31003) );
  OAI2BB1XL U16289 ( .A0N(conv_1[280]), .A1N(n29365), .B0(n29339), .Y(n35428)
         );
  OAI2BB1XL U16290 ( .A0N(conv_2[325]), .A1N(n28064), .B0(n33079), .Y(n33933)
         );
  AOI21XL U16291 ( .A0(n26714), .A1(n26709), .B0(n26710), .Y(n25447) );
  NOR2X1 U16292 ( .A(n34570), .B(n29507), .Y(n29506) );
  NOR2X1 U16293 ( .A(n30172), .B(n30924), .Y(n33811) );
  NOR2X1 U16294 ( .A(n31980), .B(n31962), .Y(n31961) );
  NOR2X1 U16295 ( .A(n33682), .B(n29455), .Y(n33195) );
  NOR2BXL U16296 ( .AN(n35301), .B(conv_1[41]), .Y(n35304) );
  AOI2BB1XL U16297 ( .A0N(conv_1[98]), .A1N(n26783), .B0(n31334), .Y(n26797)
         );
  AOI2BB1XL U16298 ( .A0N(conv_2[308]), .A1N(n29946), .B0(n35970), .Y(n35968)
         );
  AOI2BB1XL U16299 ( .A0N(conv_1[23]), .A1N(n27350), .B0(n30588), .Y(n27609)
         );
  NOR2BXL U16300 ( .AN(n36032), .B(conv_2[401]), .Y(n36034) );
  AOI2BB1XL U16301 ( .A0N(conv_1[22]), .A1N(n27338), .B0(n30588), .Y(n27350)
         );
  OR2XL U16302 ( .A(n30242), .B(n30120), .Y(n30972) );
  AOI2BB1XL U16303 ( .A0N(conv_2[502]), .A1N(n30909), .B0(n36081), .Y(n36073)
         );
  OAI2BB2XL U16304 ( .B0(n33560), .B1(n33559), .A0N(n33560), .A1N(n33559), .Y(
        n33562) );
  NOR2X1 U16305 ( .A(n27575), .B(n31363), .Y(n35453) );
  NOR2X1 U16306 ( .A(n35732), .B(n31406), .Y(n31444) );
  NOR2X1 U16307 ( .A(n34164), .B(n19194), .Y(n19198) );
  NOR2X1 U16308 ( .A(n35639), .B(n31562), .Y(n31585) );
  OAI2BB1XL U16309 ( .A0N(conv_1[10]), .A1N(n27279), .B0(n34547), .Y(n34546)
         );
  AOI2BB1XL U16310 ( .A0N(conv_2[380]), .A1N(n29444), .B0(n36025), .Y(n33415)
         );
  NOR2X1 U16311 ( .A(n34529), .B(n23079), .Y(n29445) );
  NOR2X1 U16312 ( .A(n30044), .B(n27238), .Y(n27243) );
  AOI2BB1XL U16313 ( .A0N(conv_3[95]), .A1N(n31680), .B0(n35615), .Y(n33741)
         );
  AOI2BB1XL U16314 ( .A0N(conv_2[290]), .A1N(n30888), .B0(n33135), .Y(n35955)
         );
  AOI2BB1XL U16315 ( .A0N(conv_1[366]), .A1N(n22833), .B0(n31363), .Y(n27576)
         );
  AOI32XL U16316 ( .A0(n31529), .A1(n36020), .A2(n34649), .B0(n28833), .B1(
        n33982), .Y(n28834) );
  NOR2X1 U16317 ( .A(n31137), .B(n27814), .Y(n27813) );
  NOR2X1 U16318 ( .A(n27332), .B(n27334), .Y(n26507) );
  NOR2X1 U16319 ( .A(n34626), .B(n29863), .Y(n29862) );
  NOR2X1 U16320 ( .A(n24913), .B(n27260), .Y(n27267) );
  NOR2X1 U16321 ( .A(n24913), .B(n30267), .Y(n27266) );
  AOI2BB1XL U16322 ( .A0N(conv_1[365]), .A1N(n22838), .B0(n31363), .Y(n22833)
         );
  AND2XL U16323 ( .A(n34186), .B(n31668), .Y(n31680) );
  NOR2X1 U16324 ( .A(n35957), .B(n28091), .Y(n30889) );
  NOR2X1 U16325 ( .A(n34186), .B(n31668), .Y(n31679) );
  AOI2BB1XL U16326 ( .A0N(conv_2[515]), .A1N(n27776), .B0(n28706), .Y(n33577)
         );
  NOR2X1 U16327 ( .A(n35810), .B(n19021), .Y(n26121) );
  ADDFHX2 U16328 ( .A(DP_OP_5169J1_125_4278_n39), .B(DP_OP_5169J1_125_4278_n43), .CI(n20147), .CO(n20355), .S(n20145) );
  NOR2X1 U16329 ( .A(n34292), .B(n23650), .Y(n29305) );
  OR2XL U16330 ( .A(n27273), .B(n23125), .Y(n34563) );
  NOR2X1 U16331 ( .A(n31180), .B(n31173), .Y(n31172) );
  ADDFHX2 U16332 ( .A(DP_OP_5169J1_125_4278_n44), .B(DP_OP_5169J1_125_4278_n48), .CI(n20153), .CO(n20147), .S(n20154) );
  NOR2X1 U16333 ( .A(n35515), .B(n23643), .Y(n27167) );
  AND2XL U16334 ( .A(n27237), .B(n27236), .Y(n27393) );
  AND2XL U16335 ( .A(n33580), .B(n27771), .Y(n27776) );
  NOR2X1 U16336 ( .A(n23078), .B(n23077), .Y(n29011) );
  NOR2X1 U16337 ( .A(n27451), .B(n27450), .Y(n27453) );
  ADDFX1 U16338 ( .A(conv_3[186]), .B(n32649), .CI(n32648), .CO(n31597), .S(
        n32651) );
  NOR2X1 U16339 ( .A(n35693), .B(n28798), .Y(n34245) );
  NOR2X1 U16340 ( .A(n35455), .B(n22812), .Y(n22837) );
  ADDFXL U16341 ( .A(conv_1[304]), .B(n22946), .CI(n22945), .CO(n22314), .S(
        n22947) );
  OAI21XL U16342 ( .A0(conv_1[453]), .A1(n27249), .B0(n27250), .Y(n27236) );
  NOR2X1 U16343 ( .A(n26504), .B(n26503), .Y(n27451) );
  NOR2X1 U16344 ( .A(n33770), .B(n28665), .Y(n29916) );
  OR2XL U16345 ( .A(n35884), .B(n25679), .Y(n28678) );
  NOR2X1 U16346 ( .A(intadd_1_B_2_), .B(intadd_1_n1), .Y(n35501) );
  NOR2X1 U16347 ( .A(n27554), .B(n27553), .Y(n29714) );
  NOR2X1 U16348 ( .A(n32130), .B(n31393), .Y(n31480) );
  ADDFHX2 U16349 ( .A(DP_OP_5169J1_125_4278_n49), .B(DP_OP_5169J1_125_4278_n53), .CI(n20144), .CO(n20153), .S(n20124) );
  NOR2X1 U16350 ( .A(n30267), .B(n24912), .Y(n27261) );
  AND2XL U16351 ( .A(n26131), .B(n26130), .Y(n27457) );
  AND2XL U16352 ( .A(n33953), .B(n24450), .Y(n28115) );
  AND2XL U16353 ( .A(n31134), .B(n27802), .Y(n27807) );
  NOR2X1 U16354 ( .A(n22811), .B(n22810), .Y(n30277) );
  OR2XL U16355 ( .A(n34775), .B(n25253), .Y(n26519) );
  OR2XL U16356 ( .A(n25678), .B(n25677), .Y(n34402) );
  AOI2BB1XL U16357 ( .A0N(conv_3[122]), .A1N(n30741), .B0(n30742), .Y(n35569)
         );
  NOR2X1 U16358 ( .A(n35914), .B(n28655), .Y(n29897) );
  OR2XL U16359 ( .A(n18932), .B(n18931), .Y(n34099) );
  AOI222XL U16360 ( .A0(n25808), .A1(n25807), .B0(n25808), .B1(n25806), .C0(
        n25807), .C1(n25805), .Y(n25809) );
  NAND2XL U16361 ( .A(n33058), .B(n33055), .Y(n24184) );
  ADDFX1 U16362 ( .A(DP_OP_5168J1_124_9881_n28), .B(DP_OP_5168J1_124_9881_n35), 
        .CI(n20715), .CO(n21092), .S(n20707) );
  OR2XL U16363 ( .A(n18970), .B(n18969), .Y(n25275) );
  NAND2XL U16364 ( .A(n23478), .B(n30417), .Y(n27288) );
  NAND2XL U16365 ( .A(n26500), .B(n27462), .Y(n27444) );
  ADDFXL U16366 ( .A(conv_1[318]), .B(n22438), .CI(n22437), .CO(n22950), .S(
        n22439) );
  OR2XL U16367 ( .A(n23102), .B(n23455), .Y(n23103) );
  AOI222XL U16368 ( .A0(n26977), .A1(conv_1[33]), .B0(n26977), .B1(n26976), 
        .C0(conv_1[33]), .C1(n26976), .Y(n25076) );
  AOI222XL U16369 ( .A0(pool[109]), .A1(n28362), .B0(pool[109]), .B1(n28361), 
        .C0(n28362), .C1(n28360), .Y(n28388) );
  AND2XL U16370 ( .A(n18925), .B(n18924), .Y(n30318) );
  ADDFX1 U16371 ( .A(n20688), .B(n20687), .CI(n20686), .CO(n20669), .S(n20689)
         );
  INVX1 U16372 ( .A(n26853), .Y(n31084) );
  AOI21XL U16373 ( .A0(conv_2[496]), .A1(n34232), .B0(n34233), .Y(n18925) );
  NOR4XL U16374 ( .A(n28359), .B(n28358), .C(n28379), .D(n28357), .Y(n28360)
         );
  ADDFX1 U16375 ( .A(n19709), .B(affine_2[2]), .CI(n19708), .CO(n19716), .S(
        n19712) );
  NOR2BXL U16376 ( .AN(n35849), .B(n35850), .Y(n24250) );
  OAI2BB1XL U16377 ( .A0N(conv_1[32]), .A1N(n27030), .B0(n27031), .Y(n26976)
         );
  AOI32XL U16378 ( .A0(n36056), .A1(n27427), .A2(n27426), .B0(conv_1[15]), 
        .B1(n27425), .Y(n27428) );
  INVX2 U16379 ( .A(n26853), .Y(n16645) );
  AOI2BB1XL U16380 ( .A0N(n33403), .A1N(n33429), .B0(n22217), .Y(n30461) );
  INVX1 U16381 ( .A(n31071), .Y(n32777) );
  INVX1 U16382 ( .A(n31071), .Y(n32840) );
  ADDFX1 U16383 ( .A(n20659), .B(n20658), .CI(n20657), .CO(n20666), .S(n20662)
         );
  NOR2X1 U16384 ( .A(n35858), .B(n27764), .Y(n27769) );
  NOR2X1 U16385 ( .A(n33989), .B(n27764), .Y(n23253) );
  NAND4XL U16386 ( .A(n17443), .B(n17442), .C(n17441), .D(n17440), .Y(n20634)
         );
  NOR2X1 U16387 ( .A(n25247), .B(n28948), .Y(n34292) );
  NOR2X1 U16388 ( .A(n25247), .B(n34426), .Y(n35339) );
  INVX2 U16389 ( .A(n31077), .Y(n16646) );
  NOR2X1 U16390 ( .A(n24943), .B(n36042), .Y(n24944) );
  INVX4 U16391 ( .A(n26906), .Y(n16647) );
  NOR2X1 U16392 ( .A(n24550), .B(n36042), .Y(n24551) );
  NOR2X1 U16393 ( .A(n27644), .B(n32017), .Y(n33780) );
  NOR2X1 U16394 ( .A(n29830), .B(n28948), .Y(n34344) );
  NOR2X1 U16395 ( .A(n27644), .B(n29830), .Y(n33611) );
  INVX2 U16396 ( .A(n31071), .Y(n16648) );
  NOR2X1 U16397 ( .A(n32017), .B(n34426), .Y(n33466) );
  NOR2X1 U16398 ( .A(n27644), .B(n35856), .Y(n24338) );
  NAND2XL U16399 ( .A(n27632), .B(n34444), .Y(n30051) );
  NOR2X1 U16400 ( .A(n25247), .B(n27898), .Y(n35515) );
  OAI2BB1XL U16401 ( .A0N(n33160), .A1N(n29676), .B0(n24208), .Y(n27508) );
  INVX1 U16402 ( .A(n35549), .Y(n34696) );
  NOR2X1 U16403 ( .A(n25247), .B(n28660), .Y(n35392) );
  NOR2X1 U16404 ( .A(n32017), .B(n34715), .Y(n34196) );
  NOR2X1 U16405 ( .A(n25247), .B(n28721), .Y(n30191) );
  INVX1 U16406 ( .A(n35549), .Y(n34281) );
  NOR2X1 U16407 ( .A(n35498), .B(n26717), .Y(n24316) );
  NOR2X1 U16408 ( .A(n26509), .B(n29830), .Y(n30940) );
  NOR2X1 U16409 ( .A(n35500), .B(n26717), .Y(n24318) );
  NOR2X1 U16410 ( .A(n32017), .B(n33994), .Y(n32618) );
  NOR2X1 U16411 ( .A(n29830), .B(n35499), .Y(n34211) );
  NOR2XL U16412 ( .A(n35856), .B(n35499), .Y(n32871) );
  NOR2X1 U16413 ( .A(n29830), .B(n23504), .Y(n34570) );
  INVX4 U16414 ( .A(n31384), .Y(n16649) );
  NOR2X1 U16415 ( .A(n35856), .B(n24021), .Y(n28146) );
  AOI32XL U16416 ( .A0(n17616), .A1(n17615), .A2(n17614), .B0(cursor[6]), .B1(
        n17615), .Y(n17916) );
  NOR2X1 U16417 ( .A(n35858), .B(n35499), .Y(n28132) );
  NOR2X1 U16418 ( .A(n33423), .B(n27898), .Y(n30663) );
  NOR2X1 U16419 ( .A(n25247), .B(n33994), .Y(n29364) );
  OAI2BB1XL U16420 ( .A0N(n32226), .A1N(n29676), .B0(n33442), .Y(n35641) );
  INVX1 U16421 ( .A(n35549), .Y(n34689) );
  NOR2X1 U16422 ( .A(n32017), .B(n34522), .Y(n31980) );
  NOR2X1 U16423 ( .A(n35856), .B(n26717), .Y(n23713) );
  NOR2X1 U16424 ( .A(n29830), .B(n34522), .Y(n35995) );
  NOR2X1 U16425 ( .A(n30195), .B(n32017), .Y(n33002) );
  NOR2X1 U16426 ( .A(n27848), .B(n29830), .Y(n29935) );
  AND4X2 U16427 ( .A(n22654), .B(n22653), .C(n22652), .D(n26539), .Y(n22796)
         );
  NOR2X1 U16428 ( .A(n31691), .B(n35499), .Y(n31695) );
  NOR2X1 U16429 ( .A(n35856), .B(n34522), .Y(n24302) );
  NOR2X1 U16430 ( .A(n25247), .B(n27860), .Y(n32887) );
  NOR2X1 U16431 ( .A(n35858), .B(n34522), .Y(n23867) );
  OAI2BB1XL U16432 ( .A0N(n27368), .A1N(n29676), .B0(n25246), .Y(n24536) );
  NOR2X1 U16433 ( .A(n35500), .B(n23504), .Y(n22811) );
  NOR2X1 U16434 ( .A(n32017), .B(n28721), .Y(n33480) );
  NOR2X1 U16435 ( .A(n34703), .B(n32017), .Y(n32649) );
  NOR2X1 U16436 ( .A(n33423), .B(n23504), .Y(n30058) );
  NOR2X1 U16437 ( .A(n35858), .B(n26717), .Y(n24192) );
  NOR2X1 U16438 ( .A(n25247), .B(n29136), .Y(n35404) );
  NOR2XL U16439 ( .A(n34703), .B(n18997), .Y(n23558) );
  NOR2X1 U16440 ( .A(n35500), .B(n34522), .Y(n24241) );
  NOR2X1 U16441 ( .A(n29830), .B(n29136), .Y(n32876) );
  NOR2X1 U16442 ( .A(n35498), .B(n34522), .Y(n22982) );
  NOR2X1 U16443 ( .A(n35856), .B(n27799), .Y(n27801) );
  NOR2X1 U16444 ( .A(n31691), .B(n27799), .Y(n23206) );
  NOR2X1 U16445 ( .A(n25247), .B(n26717), .Y(n35441) );
  NOR2X1 U16446 ( .A(n29830), .B(n27860), .Y(n34173) );
  INVX1 U16447 ( .A(n35549), .Y(n34682) );
  NOR2X1 U16448 ( .A(n29830), .B(n28660), .Y(n33770) );
  NOR2X1 U16449 ( .A(n29830), .B(n26717), .Y(n29526) );
  NOR2X1 U16450 ( .A(n25247), .B(n24021), .Y(n33663) );
  NOR2X1 U16451 ( .A(n30195), .B(n29830), .Y(n33620) );
  NOR2X1 U16452 ( .A(n32017), .B(n33988), .Y(n33449) );
  NOR2X1 U16453 ( .A(n25247), .B(n33988), .Y(n35296) );
  NOR2X1 U16454 ( .A(n32017), .B(n27799), .Y(n33824) );
  NOR2X1 U16455 ( .A(n25247), .B(n35499), .Y(intadd_1_B_2_) );
  INVX2 U16456 ( .A(n26853), .Y(n16650) );
  NOR2X1 U16457 ( .A(n25247), .B(n33020), .Y(n34053) );
  NOR2X1 U16458 ( .A(n29830), .B(n27799), .Y(n31137) );
  NOR2X1 U16459 ( .A(n32017), .B(n31871), .Y(n35720) );
  NOR2X1 U16460 ( .A(n27735), .B(n32017), .Y(n35831) );
  NOR2X1 U16461 ( .A(n27735), .B(n29830), .Y(n34132) );
  NOR2X1 U16462 ( .A(n35858), .B(n27799), .Y(n29739) );
  INVX1 U16463 ( .A(n35549), .Y(n34544) );
  NOR2X1 U16464 ( .A(n35498), .B(n35499), .Y(intadd_1_B_0_) );
  NOR2X2 U16465 ( .A(n27620), .B(n16654), .Y(n34742) );
  NOR2X1 U16466 ( .A(n31691), .B(n26717), .Y(n31392) );
  NOR2X1 U16467 ( .A(n25247), .B(n34715), .Y(n34557) );
  NOR2X1 U16468 ( .A(n35500), .B(n35499), .Y(intadd_1_B_1_) );
  NOR2X1 U16469 ( .A(n29830), .B(n31871), .Y(n35957) );
  NOR2X1 U16470 ( .A(n29426), .B(n26717), .Y(n26716) );
  NOR2X1 U16471 ( .A(n32017), .B(n35857), .Y(n34379) );
  INVX1 U16472 ( .A(n18856), .Y(n29675) );
  INVX1 U16473 ( .A(n18856), .Y(n24208) );
  NOR2X1 U16474 ( .A(n29830), .B(n33429), .Y(n33629) );
  NOR2X1 U16475 ( .A(n25247), .B(n33429), .Y(n29216) );
  INVX2 U16476 ( .A(n35859), .Y(n16651) );
  INVX1 U16477 ( .A(n18856), .Y(n24673) );
  INVX2 U16478 ( .A(n34461), .Y(n29136) );
  NOR2X1 U16479 ( .A(n35498), .B(n22269), .Y(n22438) );
  NOR2X1 U16480 ( .A(n35500), .B(n22269), .Y(n22949) );
  NAND2XL U16481 ( .A(n28739), .B(n33535), .Y(n29455) );
  INVX2 U16482 ( .A(n33530), .Y(n27735) );
  NAND2XL U16483 ( .A(n27632), .B(n34507), .Y(n35309) );
  AOI21XL U16484 ( .A0(n34954), .A1(n23782), .B0(n22425), .Y(n22426) );
  INVX1 U16485 ( .A(n18856), .Y(n24279) );
  NOR2X1 U16486 ( .A(n25247), .B(n19108), .Y(n28644) );
  NOR2X1 U16487 ( .A(n29830), .B(n19108), .Y(n33979) );
  AOI32XL U16488 ( .A0(n17669), .A1(n17668), .A2(n17667), .B0(cursor[6]), .B1(
        n17668), .Y(n20644) );
  NOR2X1 U16489 ( .A(n35858), .B(n22269), .Y(n23105) );
  NOR2X1 U16490 ( .A(n32017), .B(n33429), .Y(n33719) );
  AND2XL U16491 ( .A(n36020), .B(n35259), .Y(n19222) );
  NOR2X1 U16492 ( .A(n29830), .B(n28070), .Y(n36045) );
  INVX3 U16493 ( .A(n34721), .Y(n30195) );
  NOR2X1 U16494 ( .A(n32017), .B(n32016), .Y(n33699) );
  NOR2X1 U16495 ( .A(n32017), .B(n22269), .Y(n33842) );
  NOR2X1 U16496 ( .A(n31691), .B(n22269), .Y(n28756) );
  NOR2X1 U16497 ( .A(n18997), .B(n31418), .Y(n24237) );
  INVX1 U16498 ( .A(n18856), .Y(n25246) );
  NOR2X1 U16499 ( .A(n29830), .B(n32016), .Y(n34634) );
  AOI32XL U16500 ( .A0(n17911), .A1(n17910), .A2(n17909), .B0(cursor[6]), .B1(
        n17910), .Y(n20649) );
  NOR2X1 U16501 ( .A(n22269), .B(n29426), .Y(n23804) );
  NOR2X1 U16502 ( .A(n25247), .B(n35857), .Y(n27278) );
  INVX2 U16503 ( .A(n35549), .Y(n16652) );
  INVX4 U16504 ( .A(n35588), .Y(n16653) );
  BUFX2 U16505 ( .A(n17935), .Y(n19647) );
  NAND2X1 U16506 ( .A(n19037), .B(n19036), .Y(n34422) );
  INVX1 U16507 ( .A(n36042), .Y(n32181) );
  NAND3XL U16508 ( .A(n22255), .B(n22254), .C(n22253), .Y(n22256) );
  INVX1 U16509 ( .A(n36042), .Y(n32611) );
  NAND2XL U16510 ( .A(n23094), .B(n23093), .Y(n34762) );
  AOI211XL U16511 ( .A0(n35259), .A1(n19185), .B0(n19242), .C0(n19184), .Y(
        n35256) );
  AOI32X1 U16512 ( .A0(n23285), .A1(N18471), .A2(n23284), .B0(n23283), .B1(
        n28467), .Y(n34476) );
  OAI211X1 U16513 ( .A0(n23789), .A1(n26409), .B0(n23788), .C0(n23787), .Y(
        n33990) );
  INVX2 U16514 ( .A(n35336), .Y(n16654) );
  INVX1 U16515 ( .A(n26846), .Y(n26847) );
  NAND4X1 U16516 ( .A(n21106), .B(n21105), .C(n21104), .D(n21103), .Y(n34721)
         );
  INVX2 U16517 ( .A(n33912), .Y(n16655) );
  AOI21X2 U16518 ( .A0(n23055), .A1(n22153), .B0(n19201), .Y(n28070) );
  NOR2X1 U16519 ( .A(n33423), .B(n36001), .Y(n34769) );
  INVX1 U16520 ( .A(n36001), .Y(n33982) );
  NAND4X1 U16521 ( .A(n22127), .B(n22126), .C(n22125), .D(n22124), .Y(n34706)
         );
  OAI211XL U16522 ( .A0(n19143), .A1(n35135), .B0(n19142), .C0(n19141), .Y(
        n19144) );
  OAI211X1 U16523 ( .A0(n23247), .A1(n35135), .B0(n22307), .C0(n22306), .Y(
        n33535) );
  NAND3X1 U16524 ( .A(n18896), .B(n18895), .C(n18894), .Y(n33424) );
  INVX1 U16525 ( .A(n36001), .Y(n34028) );
  INVX1 U16526 ( .A(n36042), .Y(n33822) );
  AOI32X1 U16527 ( .A0(n22157), .A1(N18471), .A2(n22156), .B0(n22453), .B1(
        n28467), .Y(n34461) );
  INVX1 U16528 ( .A(n36001), .Y(n33788) );
  NAND2X1 U16529 ( .A(n19164), .B(n19163), .Y(n34450) );
  NOR2X1 U16530 ( .A(n20616), .B(n19632), .Y(n36207) );
  OAI211X1 U16531 ( .A0(N18471), .A1(n23058), .B0(n23057), .C0(n23056), .Y(
        n33530) );
  OAI211X1 U16532 ( .A0(n23247), .A1(n26575), .B0(n18772), .C0(n18771), .Y(
        n34768) );
  INVX4 U16533 ( .A(n23672), .Y(n22896) );
  OAI211X1 U16534 ( .A0(n22453), .A1(n28467), .B0(n22452), .C0(n22451), .Y(
        n34507) );
  NAND3XL U16535 ( .A(n17968), .B(n17967), .C(n17966), .Y(n17983) );
  NOR2X1 U16536 ( .A(n20618), .B(n19244), .Y(n19240) );
  OAI211X1 U16537 ( .A0(n20385), .A1(n18109), .B0(n17961), .C0(n17960), .Y(
        n17962) );
  OAI2BB1XL U16538 ( .A0N(n23274), .A1N(n22266), .B0(n22265), .Y(n22268) );
  AND2XL U16539 ( .A(n22155), .B(n22154), .Y(n22453) );
  OAI2BB1XL U16540 ( .A0N(weight_2[52]), .A1N(n18049), .B0(n18042), .Y(n18053)
         );
  OAI211XL U16541 ( .A0(N18471), .A1(n22157), .B0(n19200), .C0(n19199), .Y(
        n19201) );
  NAND3X1 U16542 ( .A(n17978), .B(n17977), .C(n17976), .Y(n24543) );
  OAI21XL U16543 ( .A0(n23282), .A1(n19106), .B0(n23058), .Y(n19107) );
  OAI211XL U16544 ( .A0(n16699), .A1(n18157), .B0(n16698), .C0(n16697), .Y(
        n20645) );
  NOR2X1 U16545 ( .A(n19244), .B(n19610), .Y(n26846) );
  INVX2 U16546 ( .A(n36042), .Y(n16657) );
  NOR2X1 U16547 ( .A(ns[1]), .B(n20615), .Y(n35227) );
  AOI211XL U16548 ( .A0(n36249), .A1(n19180), .B0(n19242), .C0(n20617), .Y(
        n35265) );
  AOI31XL U16549 ( .A0(ns[2]), .A1(n20616), .A2(n35260), .B0(n19183), .Y(
        n19184) );
  AOI2BB2XL U16550 ( .B0(n23017), .B1(n22448), .A0N(N18471), .A1N(n22265), .Y(
        n18894) );
  NAND2XL U16551 ( .A(n19121), .B(n19120), .Y(n22267) );
  OAI211XL U16552 ( .A0(n22401), .A1(n19181), .B0(n19035), .C0(n19034), .Y(
        n23092) );
  INVX2 U16553 ( .A(n36056), .Y(n16658) );
  OAI211XL U16554 ( .A0(n16854), .A1(n18157), .B0(n16853), .C0(n16852), .Y(
        n17918) );
  OAI211XL U16555 ( .A0(n16986), .A1(n18157), .B0(n16985), .C0(n16984), .Y(
        n20646) );
  OAI211XL U16556 ( .A0(n17041), .A1(n18157), .B0(n17040), .C0(n17039), .Y(
        n33554) );
  NAND2XL U16557 ( .A(n18947), .B(n18946), .Y(n22123) );
  AND2X1 U16558 ( .A(n18739), .B(n18738), .Y(n23247) );
  AND2XL U16559 ( .A(n18943), .B(n18942), .Y(n22807) );
  AOI222XL U16560 ( .A0(n23782), .A1(n23278), .B0(n23277), .B1(n23276), .C0(
        n23781), .C1(n23272), .Y(n23058) );
  OAI211XL U16561 ( .A0(n23789), .A1(n19106), .B0(n19105), .C0(n19104), .Y(
        n22422) );
  NAND2XL U16562 ( .A(n21099), .B(n21098), .Y(n22848) );
  AND4X2 U16563 ( .A(n19072), .B(n19071), .C(n19070), .D(n19069), .Y(n23282)
         );
  AOI22XL U16564 ( .A0(n28414), .A1(n22212), .B0(n28556), .B1(n22843), .Y(
        n21106) );
  NOR2X1 U16565 ( .A(N18471), .B(n19226), .Y(n19187) );
  OAI211XL U16566 ( .A0(n17009), .A1(n18157), .B0(n17008), .C0(n17007), .Y(
        n20648) );
  AND2X1 U16567 ( .A(n20617), .B(ns[1]), .Y(n19183) );
  INVX2 U16568 ( .A(n21731), .Y(n21749) );
  NAND2XL U16569 ( .A(n18789), .B(n18788), .Y(n22204) );
  OAI2BB1X2 U16570 ( .A0N(n18184), .A1N(n18183), .B0(n19180), .Y(ns[1]) );
  NOR2X1 U16571 ( .A(ns[2]), .B(n19244), .Y(n20617) );
  NAND2XL U16572 ( .A(n18787), .B(n18786), .Y(n22211) );
  INVX2 U16573 ( .A(n28479), .Y(n16659) );
  INVX1 U16574 ( .A(n19185), .Y(ns[2]) );
  INVX2 U16575 ( .A(n35198), .Y(n16660) );
  BUFX3 U16576 ( .A(n18845), .Y(n27429) );
  INVX1 U16577 ( .A(n28739), .Y(n29830) );
  INVX1 U16578 ( .A(n27632), .Y(n25247) );
  NOR2X1 U16579 ( .A(n22550), .B(n26621), .Y(n17812) );
  NOR2X1 U16580 ( .A(n22717), .B(n18782), .Y(n17809) );
  INVX1 U16581 ( .A(n31924), .Y(n32017) );
  NAND4BXL U16582 ( .AN(n18985), .B(n18984), .C(n18983), .D(n18982), .Y(n24467) );
  NOR2X1 U16583 ( .A(n18321), .B(n29178), .Y(n18292) );
  NOR2X1 U16584 ( .A(n18321), .B(n32135), .Y(n18666) );
  BUFX4 U16585 ( .A(n16703), .Y(n19475) );
  NOR2X1 U16586 ( .A(n18321), .B(n29932), .Y(n20874) );
  NOR2X1 U16587 ( .A(cs[1]), .B(n18167), .Y(n18163) );
  BUFX4 U16588 ( .A(n16709), .Y(n19097) );
  NAND4BXL U16589 ( .AN(n18980), .B(n18979), .C(n18978), .D(n18977), .Y(n31924) );
  NOR2X1 U16590 ( .A(n22759), .B(n26039), .Y(n35255) );
  INVX2 U16591 ( .A(n26263), .Y(n16661) );
  NOR2X1 U16592 ( .A(n18321), .B(n29655), .Y(n18611) );
  NOR2X1 U16593 ( .A(n22716), .B(n35239), .Y(n17864) );
  NOR2X1 U16594 ( .A(n16715), .B(n35239), .Y(n17788) );
  NOR2X1 U16595 ( .A(n16715), .B(n26279), .Y(n17888) );
  NOR2X1 U16596 ( .A(n22716), .B(n26279), .Y(n17899) );
  OAI31X1 U16597 ( .A0(in_valid_1), .A1(n18179), .A2(n18189), .B0(n18178), .Y(
        n18180) );
  NAND4BXL U16598 ( .AN(n18906), .B(n18905), .C(n18904), .D(n18903), .Y(n29046) );
  INVX4 U16599 ( .A(n22740), .Y(n16662) );
  NAND4BXL U16600 ( .AN(n18901), .B(n18900), .C(n18899), .D(n18898), .Y(n28739) );
  NAND2X2 U16601 ( .A(n22759), .B(n28290), .Y(n18116) );
  NOR2X1 U16602 ( .A(n22765), .B(n26285), .Y(n21751) );
  INVX2 U16603 ( .A(n28349), .Y(n16663) );
  OAI21X1 U16604 ( .A0(cs[3]), .A1(n18188), .B0(n18187), .Y(n19244) );
  OAI2BB1XL U16605 ( .A0N(n19008), .A1N(filter_1[47]), .B0(n18725), .Y(n18729)
         );
  NOR2X1 U16606 ( .A(n16715), .B(n29958), .Y(n20763) );
  INVX2 U16607 ( .A(n35200), .Y(n16664) );
  INVX16 U16608 ( .A(n18239), .Y(n22759) );
  INVX2 U16609 ( .A(n28553), .Y(n16665) );
  INVX2 U16610 ( .A(n22369), .Y(n18815) );
  INVX3 U16611 ( .A(n18776), .Y(n16666) );
  NOR2X1 U16612 ( .A(n18173), .B(n19227), .Y(n18184) );
  INVX2 U16613 ( .A(n28577), .Y(n16667) );
  NOR2X1 U16614 ( .A(n16715), .B(n30124), .Y(n20845) );
  NOR2X1 U16615 ( .A(n16715), .B(n31678), .Y(n18532) );
  INVX2 U16616 ( .A(n22616), .Y(n16668) );
  OAI2BB1XL U16617 ( .A0N(n20605), .A1N(filter_2[5]), .B0(n18897), .Y(n18901)
         );
  NOR2X1 U16618 ( .A(counter[4]), .B(n17017), .Y(n17010) );
  NOR2X1 U16619 ( .A(n18160), .B(n18177), .Y(n18190) );
  NOR2X1 U16620 ( .A(n20432), .B(n21358), .Y(n21167) );
  NOR2X1 U16621 ( .A(n20473), .B(n21358), .Y(n21319) );
  INVX2 U16622 ( .A(n26474), .Y(n16671) );
  NOR2X1 U16623 ( .A(n36246), .B(n19470), .Y(n21173) );
  NOR2X1 U16624 ( .A(n22226), .B(n21358), .Y(n21114) );
  NOR2X1 U16625 ( .A(n22716), .B(n33469), .Y(n19426) );
  NOR2X1 U16626 ( .A(n36246), .B(n21147), .Y(n20442) );
  NOR2X1 U16627 ( .A(n36246), .B(n21295), .Y(n21296) );
  NOR2X1 U16628 ( .A(n36246), .B(n19558), .Y(n20562) );
  NOR2X1 U16629 ( .A(n22716), .B(n32175), .Y(n19528) );
  NOR2X1 U16630 ( .A(n28292), .B(n16701), .Y(n34984) );
  NOR2X1 U16631 ( .A(n22716), .B(n31864), .Y(n19560) );
  NOR2X1 U16632 ( .A(n22716), .B(n32793), .Y(n19546) );
  NOR2X1 U16633 ( .A(n20514), .B(n21358), .Y(n21329) );
  NOR2X1 U16634 ( .A(n36246), .B(n22489), .Y(n21639) );
  NOR2X1 U16635 ( .A(n36246), .B(n24043), .Y(n20742) );
  NOR2X1 U16636 ( .A(n24042), .B(n21358), .Y(n34904) );
  OAI2BB1XL U16637 ( .A0N(n20605), .A1N(filter_3[5]), .B0(n18976), .Y(n18980)
         );
  INVX2 U16638 ( .A(n18463), .Y(n16672) );
  NOR2X1 U16639 ( .A(n20164), .B(n18172), .Y(n18773) );
  NOR2X1 U16640 ( .A(n19245), .B(n18170), .Y(n20358) );
  NOR2X1 U16641 ( .A(n36246), .B(n22683), .Y(n19834) );
  NOR2X1 U16642 ( .A(n19181), .B(n16701), .Y(n28556) );
  NOR2X1 U16643 ( .A(n18185), .B(n18186), .Y(n18182) );
  NOR2X1 U16644 ( .A(n36246), .B(n22745), .Y(n21768) );
  NOR2X1 U16645 ( .A(n22716), .B(n30233), .Y(n21067) );
  NOR2X1 U16646 ( .A(n36246), .B(n20803), .Y(n25977) );
  NOR2X1 U16647 ( .A(n36246), .B(n25936), .Y(n21863) );
  NOR2X1 U16648 ( .A(n20601), .B(n17028), .Y(n17011) );
  NOR2X1 U16649 ( .A(n36246), .B(n21858), .Y(n25939) );
  NOR2X1 U16650 ( .A(n22488), .B(n21358), .Y(n21643) );
  NOR2X1 U16651 ( .A(n20601), .B(n17029), .Y(n18159) );
  NOR2X1 U16652 ( .A(n20600), .B(n20599), .Y(n20602) );
  AOI2BB1XL U16653 ( .A0N(counter[2]), .A1N(counter[1]), .B0(n20601), .Y(
        n20604) );
  NOR2X1 U16654 ( .A(n16721), .B(n16701), .Y(n23783) );
  INVX8 U16655 ( .A(n22716), .Y(n16673) );
  INVX4 U16656 ( .A(n16701), .Y(n34827) );
  NOR2X1 U16657 ( .A(n18156), .B(n18158), .Y(n18191) );
  NOR2X1 U16658 ( .A(n20164), .B(n20163), .Y(n36122) );
  NAND2XL U16659 ( .A(counter[3]), .B(n20600), .Y(n20601) );
  NAND2X1 U16660 ( .A(cs[3]), .B(n18160), .Y(n18187) );
  AOI221X1 U16661 ( .A0(in_valid_1), .A1(n18161), .B0(n18179), .B1(cs[1]), 
        .C0(cs[2]), .Y(n18162) );
  INVX1 U16662 ( .A(counter[4]), .Y(n20600) );
  INVX1 U16663 ( .A(counter[2]), .Y(n19246) );
  INVX1 U16664 ( .A(counter[3]), .Y(n19247) );
  NOR2X1 U16665 ( .A(cs[1]), .B(cs[2]), .Y(n18160) );
  NOR2X1 U16666 ( .A(counter[6]), .B(counter[5]), .Y(n20165) );
  INVX4 U16667 ( .A(in_valid_2), .Y(n18179) );
  NOR2X1 U16668 ( .A(n33416), .B(n36025), .Y(n36023) );
  OAI211XL U16669 ( .A0(n34789), .A1(n28160), .B0(n34669), .C0(n28159), .Y(
        n14944) );
  AOI22XL U16670 ( .A0(conv_2[388]), .A1(n28156), .B0(n28155), .B1(n28154), 
        .Y(n28158) );
  NOR2X1 U16671 ( .A(n36245), .B(n23052), .Y(n18535) );
  OAI211XL U16672 ( .A0(n33442), .A1(n33134), .B0(n34281), .C0(n33133), .Y(
        n16089) );
  AOI22XL U16673 ( .A0(conv_1[373]), .A1(n33130), .B0(n33129), .B1(n33128), 
        .Y(n33132) );
  NAND4BX2 U16674 ( .AN(n18839), .B(n18838), .C(n18837), .D(n18836), .Y(n30672) );
  INVX2 U16675 ( .A(n22105), .Y(n36100) );
  ADDFHX1 U16676 ( .A(DP_OP_5170J1_126_4278_n25), .B(n28400), .CI(n28399), 
        .CO(n33342), .S(n24565) );
  NAND2X1 U16677 ( .A(n19098), .B(n19221), .Y(n18119) );
  OAI211X1 U16678 ( .A0(n34520), .A1(n32204), .B0(n16649), .C0(n32203), .Y(
        n15484) );
  NAND2XL U16679 ( .A(n33351), .B(n33350), .Y(n16530) );
  NAND2X4 U16680 ( .A(n20735), .B(n17923), .Y(n18043) );
  NOR2X1 U16681 ( .A(n19221), .B(n21830), .Y(n17923) );
  INVX1 U16682 ( .A(n17962), .Y(n19638) );
  ADDFHX1 U16683 ( .A(DP_OP_5169J1_125_4278_n25), .B(n28213), .CI(n28212), 
        .CO(n33332), .S(n24548) );
  AOI2BB1XL U16684 ( .A0N(conv_2[83]), .A1N(n35874), .B0(n30924), .Y(n28744)
         );
  AOI2BB1XL U16685 ( .A0N(conv_2[82]), .A1N(n30166), .B0(n30924), .Y(n35874)
         );
  OAI211XL U16686 ( .A0(n34676), .A1(n32677), .B0(n33815), .C0(n32676), .Y(
        n15144) );
  OAI211XL U16687 ( .A0(conv_2[89]), .A1(n32675), .B0(n33982), .C0(n32674), 
        .Y(n32676) );
  AOI22XL U16688 ( .A0(conv_2[88]), .A1(n32673), .B0(n32672), .B1(n32671), .Y(
        n32675) );
  ADDFHX1 U16689 ( .A(DP_OP_5166J1_122_9881_n21), .B(DP_OP_5166J1_122_9881_n17), .CI(n25068), .CO(n33405), .S(n22119) );
  ADDFHX1 U16690 ( .A(DP_OP_5166J1_122_9881_n16), .B(DP_OP_5166J1_122_9881_n14), .CI(n33405), .CO(n33406), .S(n25070) );
  OR2X1 U16691 ( .A(n19902), .B(n34981), .Y(n21710) );
  NOR2X2 U16692 ( .A(n33989), .B(n16654), .Y(n34581) );
  NAND2XL U16693 ( .A(n33369), .B(n33368), .Y(n16564) );
  AOI22XL U16694 ( .A0(affine_2[15]), .A1(n33367), .B0(n16674), .B1(n33366), 
        .Y(n33369) );
  NOR2X1 U16695 ( .A(n35269), .B(n21358), .Y(n16725) );
  INVX8 U16696 ( .A(n19855), .Y(n35269) );
  INVX4 U16697 ( .A(N17631), .Y(n19855) );
  CLKINVX2 U16698 ( .A(n24572), .Y(n28611) );
  NAND2XL U16699 ( .A(conv_3[269]), .B(n33909), .Y(n33908) );
  AOI22XL U16700 ( .A0(conv_3[268]), .A1(n33907), .B0(n33906), .B1(n33905), 
        .Y(n33909) );
  AOI222X1 U16701 ( .A0(n28723), .A1(n28722), .B0(n28723), .B1(conv_3[259]), 
        .C0(n28722), .C1(conv_3[259]), .Y(n28724) );
  AOI2BB1X2 U16702 ( .A0N(conv_3[258]), .A1N(n29414), .B0(n29415), .Y(n28722)
         );
  AND2X2 U16703 ( .A(n28292), .B(n36244), .Y(n28407) );
  OR2X2 U16704 ( .A(n35599), .B(n35600), .Y(n35601) );
  OAI211X1 U16705 ( .A0(n34789), .A1(n32168), .B0(n16649), .C0(n32167), .Y(
        n15694) );
  ADDFHX1 U16706 ( .A(DP_OP_5166J1_122_9881_n28), .B(DP_OP_5166J1_122_9881_n35), .CI(n20709), .CO(n22118), .S(n20710) );
  OAI211XL U16707 ( .A0(conv_3[14]), .A1(n33158), .B0(n33157), .C0(n33156), 
        .Y(n33159) );
  AOI22XL U16708 ( .A0(conv_3[13]), .A1(n33155), .B0(n33154), .B1(n33153), .Y(
        n33158) );
  ADDFHX1 U16709 ( .A(conv_3[7]), .B(n34379), .CI(n24376), .CO(n31194), .S(
        n24377) );
  OAI2BB2XL U16710 ( .B0(n24371), .B1(n32996), .A0N(conv_3[6]), .A1N(n31427), 
        .Y(n24376) );
  INVXL U16711 ( .A(n31026), .Y(n23752) );
  XOR2X1 U16712 ( .A(affine_2[31]), .B(n33345), .Y(n33348) );
  AOI22XL U16713 ( .A0(affine_2[31]), .A1(n33367), .B0(n16674), .B1(n33349), 
        .Y(n33351) );
  OAI2BB1X2 U16714 ( .A0N(weight_2[49]), .A1N(n18049), .B0(n18015), .Y(n19626)
         );
  NOR4X1 U16715 ( .A(n18014), .B(n18013), .C(n18012), .D(n18011), .Y(n18015)
         );
  MXI2X1 U16716 ( .A(n19629), .B(n19626), .S0(n19611), .Y(n19612) );
  INVX2 U16717 ( .A(n19626), .Y(n19629) );
  NAND2XL U16718 ( .A(n33341), .B(n33340), .Y(n16546) );
  ADDFHX1 U16719 ( .A(DP_OP_5169J1_125_4278_n54), .B(DP_OP_5169J1_125_4278_n58), .CI(n20156), .CO(n20144), .S(n20157) );
  AOI22XL U16720 ( .A0(n33563), .A1(n33411), .B0(affine_1[29]), .B1(n33561), 
        .Y(n33413) );
  NAND2XL U16721 ( .A(n33413), .B(n33412), .Y(n16492) );
  NOR2X4 U16722 ( .A(n36245), .B(n18750), .Y(n21887) );
  NAND2X4 U16723 ( .A(n22896), .B(filter_2_bias[5]), .Y(n35859) );
  AOI22XL U16724 ( .A0(n33563), .A1(n33076), .B0(affine_1[9]), .B1(n33561), 
        .Y(n33078) );
  AOI2BB1XL U16725 ( .A0N(conv_3[125]), .A1N(n31398), .B0(n31399), .Y(n32662)
         );
  AOI21XL U16726 ( .A0(conv_3[121]), .A1(n27514), .B0(n27513), .Y(n23686) );
  NOR2X1 U16727 ( .A(n36245), .B(n16715), .Y(n16706) );
  NAND2XL U16728 ( .A(n23276), .B(n23784), .Y(n19104) );
  NAND2XL U16729 ( .A(conv_3[134]), .B(n34786), .Y(n34785) );
  AOI222XL U16730 ( .A0(n35570), .A1(n35569), .B0(n35570), .B1(conv_3[123]), 
        .C0(n35569), .C1(conv_3[123]), .Y(n23688) );
  OAI32XL U16731 ( .A0(conv_3[133]), .A1(n34784), .A2(n34783), .B0(n34782), 
        .B1(n34781), .Y(n34786) );
  NAND2XL U16732 ( .A(n34784), .B(n34783), .Y(n34782) );
  AND2X2 U16733 ( .A(filter_1_bias[5]), .B(n22896), .Y(n35549) );
  OR2XL U16734 ( .A(n35549), .B(n33255), .Y(n16420) );
  OAI22XL U16735 ( .A0(n16654), .A1(n33254), .B0(n35302), .B1(n33253), .Y(
        n33255) );
  AOI2BB1XL U16736 ( .A0N(conv_1[37]), .A1N(n35287), .B0(n35289), .Y(n27300)
         );
  AOI2BB1XL U16737 ( .A0N(conv_1[36]), .A1N(n35281), .B0(n35289), .Y(n35287)
         );
  OAI2BB2XL U16738 ( .B0(conv_1[43]), .B1(n33252), .A0N(conv_1[43]), .A1N(
        n33252), .Y(n33254) );
  NOR2X2 U16739 ( .A(n19246), .B(n16675), .Y(n16676) );
  INVX1 U16740 ( .A(n18003), .Y(n19640) );
  AOI22XL U16741 ( .A0(affine_2[47]), .A1(n33367), .B0(n16674), .B1(n33339), 
        .Y(n33341) );
  MXI2X2 U16742 ( .A(n19650), .B(n19647), .S0(n19636), .Y(n19637) );
  INVX3 U16743 ( .A(n19647), .Y(n19650) );
  NAND2XL U16744 ( .A(counter[1]), .B(n36248), .Y(n16675) );
  NAND2X1 U16745 ( .A(n17988), .B(n19246), .Y(n17029) );
  INVX2 U16746 ( .A(n26376), .Y(n26274) );
  AOI22XL U16747 ( .A0(n22362), .A1(n22121), .B0(n22369), .B1(n22122), .Y(
        n18942) );
  AOI22XL U16748 ( .A0(n22370), .A1(n22171), .B0(n21100), .B1(n22170), .Y(
        n18943) );
  OAI21XL U16749 ( .A0(n19098), .A1(n19221), .B0(n18119), .Y(n18049) );
  NAND4BX1 U16750 ( .AN(n18930), .B(n18929), .C(n18928), .D(n18927), .Y(n28068) );
  AOI22XL U16751 ( .A0(n19007), .A1(filter_2[27]), .B0(n19005), .B1(
        filter_2[15]), .Y(n18929) );
  AOI22XL U16752 ( .A0(n19004), .A1(filter_2[33]), .B0(n16676), .B1(
        filter_2[39]), .Y(n18928) );
  INVXL U16753 ( .A(n26262), .Y(n26279) );
  AOI22XL U16754 ( .A0(n34963), .A1(n35061), .B0(n26451), .B1(n35054), .Y(
        n24826) );
  AOI22XL U16755 ( .A0(pixel[52]), .A1(n22021), .B0(pixel[57]), .B1(n19098), 
        .Y(n19069) );
  NAND2XL U16756 ( .A(n18756), .B(n18755), .Y(n23242) );
  NAND2XL U16757 ( .A(n18754), .B(n18753), .Y(n23243) );
  NAND2XL U16758 ( .A(n18752), .B(n18751), .Y(n23241) );
  NOR2XL U16759 ( .A(N18014), .B(n36244), .Y(n23278) );
  NOR2XL U16760 ( .A(N18014), .B(n16721), .Y(n23272) );
  OAI21XL U16761 ( .A0(n28292), .A1(n25109), .B0(n18350), .Y(n24707) );
  NAND2XL U16762 ( .A(n23055), .B(n19099), .Y(n26085) );
  AOI211XL U16763 ( .A0(n22770), .A1(conv_3[78]), .B0(n18611), .C0(n18610), 
        .Y(n35126) );
  INVXL U16764 ( .A(n28068), .Y(n35856) );
  NAND4BX1 U16765 ( .AN(n18923), .B(n18922), .C(n18921), .D(n18920), .Y(n28128) );
  AOI22XL U16766 ( .A0(n19008), .A1(filter_2[44]), .B0(n19005), .B1(
        filter_2[14]), .Y(n18922) );
  AOI22XL U16767 ( .A0(n19006), .A1(filter_2[8]), .B0(n19004), .B1(
        filter_2[32]), .Y(n18920) );
  AOI22XL U16768 ( .A0(n19007), .A1(filter_2[26]), .B0(n16676), .B1(
        filter_2[38]), .Y(n18921) );
  NAND2XL U16769 ( .A(n18960), .B(n18959), .Y(n22305) );
  AOI22XL U16770 ( .A0(n22362), .A1(n19050), .B0(n22369), .B1(n22802), .Y(
        n18960) );
  NAND2XL U16771 ( .A(n18763), .B(n18762), .Y(n19052) );
  AOI22XL U16772 ( .A0(n16716), .A1(pixel[2]), .B0(n25299), .B1(pixel[0]), .Y(
        n18762) );
  NOR2X2 U16773 ( .A(n18815), .B(n35241), .Y(n26376) );
  NAND2XL U16774 ( .A(n18759), .B(n18758), .Y(n23244) );
  NOR2X2 U16775 ( .A(n19181), .B(n35241), .Y(n26262) );
  NAND2XL U16776 ( .A(n18749), .B(n18748), .Y(n23249) );
  AOI22XL U16777 ( .A0(n22362), .A1(n22802), .B0(n22369), .B1(n19050), .Y(
        n18749) );
  NOR2X1 U16778 ( .A(n36244), .B(n19221), .Y(n23274) );
  NAND2XL U16779 ( .A(n18731), .B(n18730), .Y(n22171) );
  INVXL U16780 ( .A(n22844), .Y(n22401) );
  INVXL U16781 ( .A(n17866), .Y(n17143) );
  INVXL U16782 ( .A(n17821), .Y(n17188) );
  AOI22XL U16783 ( .A0(n25306), .A1(conv_1[140]), .B0(n16662), .B1(conv_1[155]), .Y(n22581) );
  AOI22XL U16784 ( .A0(n25306), .A1(conv_1[86]), .B0(n16673), .B1(conv_1[116]), 
        .Y(n22602) );
  AOI2BB2XL U16785 ( .B0(n36245), .B1(n28500), .A0N(n28499), .A1N(n36245), .Y(
        n26593) );
  AOI22XL U16786 ( .A0(n25306), .A1(conv_1[146]), .B0(n16662), .B1(conv_1[161]), .Y(n22598) );
  AOI22XL U16787 ( .A0(n34963), .A1(n25531), .B0(n26276), .B1(n25533), .Y(
        n24985) );
  AOI211XL U16788 ( .A0(conv_2[5]), .A1(n22759), .B0(n18238), .C0(n18237), .Y(
        n25518) );
  AOI22XL U16789 ( .A0(n16662), .A1(conv_3[37]), .B0(n22615), .B1(conv_3[52]), 
        .Y(n18524) );
  NOR4XL U16790 ( .A(n18035), .B(n18034), .C(n18033), .D(n18032), .Y(n18036)
         );
  OAI211XL U16791 ( .A0(n20365), .A1(n18127), .B0(n18126), .C0(n18125), .Y(
        n18128) );
  OAI211XL U16792 ( .A0(n20371), .A1(n18121), .B0(n18114), .C0(n18113), .Y(
        n18132) );
  INVXL U16793 ( .A(n18128), .Y(n24571) );
  OAI2BB1X1 U16794 ( .A0N(weight_2[53]), .A1N(n18049), .B0(n18048), .Y(n24560)
         );
  MXI2XL U16795 ( .A(n19613), .B(n19614), .S0(n18053), .Y(n24562) );
  INVXL U16796 ( .A(n24560), .Y(n24561) );
  NAND2X1 U16797 ( .A(n19228), .B(n19246), .Y(n17027) );
  AOI22XL U16798 ( .A0(n25306), .A1(conv_1[288]), .B0(n16662), .B1(conv_1[303]), .Y(n19800) );
  AOI22XL U16799 ( .A0(n25306), .A1(conv_1[348]), .B0(n16662), .B1(conv_1[363]), .Y(n19796) );
  INVXL U16800 ( .A(n21959), .Y(n21998) );
  NAND4BXL U16801 ( .AN(n18829), .B(n18828), .C(n18827), .D(n18826), .Y(n27231) );
  AOI22XL U16802 ( .A0(n19009), .A1(filter_1[21]), .B0(n19007), .B1(
        filter_1[27]), .Y(n18827) );
  INVXL U16803 ( .A(n22015), .Y(n21953) );
  NAND4BX1 U16804 ( .AN(n18990), .B(n18989), .C(n18988), .D(n18987), .Y(n29677) );
  AOI22XL U16805 ( .A0(n19009), .A1(filter_3[21]), .B0(n19006), .B1(
        filter_3[9]), .Y(n18988) );
  AOI22XL U16806 ( .A0(n19007), .A1(filter_3[27]), .B0(n19005), .B1(
        filter_3[15]), .Y(n18987) );
  AOI22XL U16807 ( .A0(n19004), .A1(filter_3[33]), .B0(n16676), .B1(
        filter_3[39]), .Y(n18989) );
  AOI22XL U16808 ( .A0(n34963), .A1(n28437), .B0(n28436), .B1(n28372), .Y(
        n26608) );
  AOI22XL U16809 ( .A0(n25306), .A1(conv_1[89]), .B0(n16662), .B1(conv_1[104]), 
        .Y(n22715) );
  NAND4BXL U16810 ( .AN(n18824), .B(n18823), .C(n18822), .D(n18821), .Y(n27230) );
  NAND2XL U16811 ( .A(N18471), .B(n16721), .Y(n20755) );
  NOR2X1 U16812 ( .A(n20818), .B(n20817), .Y(n21035) );
  INVXL U16813 ( .A(n19097), .Y(n20726) );
  AOI22XL U16814 ( .A0(n36244), .A1(n25560), .B0(n34963), .B1(n25558), .Y(
        n25015) );
  AOI22XL U16815 ( .A0(n34963), .A1(n25588), .B0(n34984), .B1(n24747), .Y(
        n24073) );
  NAND2XL U16816 ( .A(n22616), .B(n26263), .Y(n22030) );
  INVX2 U16817 ( .A(n16723), .Y(n18750) );
  AOI22XL U16818 ( .A0(n34963), .A1(n28371), .B0(n26262), .B1(n26261), .Y(
        n26266) );
  NOR4BBXL U16819 ( .AN(n27067), .BN(n26236), .C(n26272), .D(n26271), .Y(
        n26255) );
  AOI22XL U16820 ( .A0(n22690), .A1(conv_3[194]), .B0(n22615), .B1(conv_3[239]), .Y(n18654) );
  INVXL U16821 ( .A(n18475), .Y(n18782) );
  NAND2XL U16822 ( .A(n18765), .B(n18764), .Y(n19051) );
  AOI22XL U16823 ( .A0(pixel[53]), .A1(n22021), .B0(pixel[51]), .B1(n21954), 
        .Y(n18869) );
  INVX2 U16824 ( .A(n17029), .Y(n19006) );
  AOI22XL U16825 ( .A0(pixel[44]), .A1(n22021), .B0(pixel[43]), .B1(n16734), 
        .Y(n19076) );
  INVXL U16826 ( .A(n22889), .Y(n21095) );
  OR2X1 U16827 ( .A(n20164), .B(counter[2]), .Y(n18157) );
  NAND2XL U16828 ( .A(ns[2]), .B(ns[0]), .Y(n20615) );
  INVXL U16829 ( .A(n24562), .Y(n28398) );
  NOR2X2 U16830 ( .A(counter[3]), .B(n17027), .Y(n20605) );
  AOI21XL U16831 ( .A0(n25399), .A1(n25398), .B0(n25397), .Y(n25401) );
  AOI22XL U16832 ( .A0(n36245), .A1(n24624), .B0(n25396), .B1(n26374), .Y(
        n26554) );
  NAND2XL U16833 ( .A(n25117), .B(n25484), .Y(n25481) );
  NOR2X1 U16834 ( .A(n26555), .B(n25123), .Y(n22672) );
  NOR2X1 U16835 ( .A(n23419), .B(n24943), .Y(n23420) );
  NOR2X1 U16836 ( .A(n23417), .B(n33421), .Y(n23419) );
  NOR2X1 U16837 ( .A(n25120), .B(n25123), .Y(n25121) );
  AOI211XL U16838 ( .A0(n21100), .A1(n25127), .B0(n25126), .C0(n25125), .Y(
        n25493) );
  NOR2X1 U16839 ( .A(n25124), .B(n25123), .Y(n25126) );
  AOI211XL U16840 ( .A0(n25399), .A1(n25488), .B0(n24965), .C0(n24964), .Y(
        n25128) );
  INVXL U16841 ( .A(n24715), .Y(n25120) );
  NAND2X1 U16842 ( .A(n28290), .B(n26172), .Y(n28277) );
  OAI2BB1XL U16843 ( .A0N(n28289), .A1N(n25380), .B0(n25379), .Y(n28427) );
  AOI211XL U16844 ( .A0(n25399), .A1(n25378), .B0(n26382), .C0(n25377), .Y(
        n25379) );
  AOI22XL U16845 ( .A0(n25299), .A1(conv_2[33]), .B0(n22615), .B1(conv_2[78]), 
        .Y(n20958) );
  NOR2X1 U16846 ( .A(n35195), .B(n34954), .Y(n19767) );
  NOR2X1 U16847 ( .A(n23097), .B(n24486), .Y(n29878) );
  NOR2X1 U16848 ( .A(n22899), .B(n24555), .Y(n34614) );
  AOI22XL U16849 ( .A0(n28528), .A1(n26570), .B0(n34963), .B1(n26569), .Y(
        n26408) );
  INVXL U16850 ( .A(n27231), .Y(n35498) );
  INVXL U16851 ( .A(n34984), .Y(n26473) );
  INVXL U16852 ( .A(n19767), .Y(n24056) );
  AOI22XL U16853 ( .A0(n18658), .A1(conv_3[124]), .B0(n22615), .B1(conv_3[169]), .Y(n18490) );
  INVXL U16854 ( .A(n29677), .Y(n29426) );
  NOR4XL U16855 ( .A(n25422), .B(n25421), .C(n25420), .D(n25419), .Y(n25427)
         );
  AOI2BB2XL U16856 ( .B0(pool[4]), .B1(n25411), .A0N(n25410), .A1N(n25409), 
        .Y(n25432) );
  AOI22XL U16857 ( .A0(n34963), .A1(n34846), .B0(n16671), .B1(n26532), .Y(
        n26375) );
  AOI2BB2XL U16858 ( .B0(n36245), .B1(n28411), .A0N(n28416), .A1N(n36245), .Y(
        n26639) );
  OAI2BB1XL U16859 ( .A0N(conv_1[516]), .A1N(n27267), .B0(n30267), .Y(n25258)
         );
  AOI2BB1XL U16860 ( .A0N(conv_1[489]), .A1N(n29982), .B0(n35534), .Y(n29992)
         );
  AOI2BB1XL U16861 ( .A0N(conv_1[394]), .A1N(n30759), .B0(n30760), .Y(n27637)
         );
  INVXL U16862 ( .A(n27230), .Y(n35500) );
  AOI22XL U16863 ( .A0(n22847), .A1(n22846), .B0(n16659), .B1(n22845), .Y(
        n22853) );
  AOI222XL U16864 ( .A0(n26116), .A1(n26057), .B0(n26116), .B1(n26056), .C0(
        n26057), .C1(n26055), .Y(n26110) );
  NOR4BXL U16865 ( .AN(n26054), .B(n26115), .C(n26053), .D(n26052), .Y(n26055)
         );
  AOI22XL U16866 ( .A0(n36245), .A1(n25618), .B0(n25621), .B1(n28292), .Y(
        n24783) );
  OAI2BB2XL U16867 ( .B0(n18405), .B1(n18404), .A0N(pool[89]), .A1N(n18403), 
        .Y(n18448) );
  INVXL U16868 ( .A(n34132), .Y(n34130) );
  AOI2BB1XL U16869 ( .A0N(conv_2[368]), .A1N(n29507), .B0(n27273), .Y(n29492)
         );
  INVXL U16870 ( .A(n34570), .Y(n27273) );
  AOI222XL U16871 ( .A0(conv_2[349]), .A1(n24192), .B0(conv_2[349]), .B1(
        n24193), .C0(n24192), .C1(n24193), .Y(n33924) );
  AOI222XL U16872 ( .A0(n29062), .A1(n29063), .B0(n29062), .B1(conv_2[274]), 
        .C0(n29063), .C1(conv_2[274]), .Y(n18955) );
  AOI2BB1XL U16873 ( .A0N(n30075), .A1N(n30071), .B0(n34344), .Y(n34351) );
  MXI2X1 U16874 ( .A(n22378), .B(n22377), .S0(N18471), .Y(n27691) );
  OAI32XL U16875 ( .A0(n19221), .A1(n22346), .A2(n22345), .B0(N18014), .B1(
        n22344), .Y(n22378) );
  OAI32XL U16876 ( .A0(n19221), .A1(n22376), .A2(n22375), .B0(N18014), .B1(
        n22374), .Y(n22377) );
  AOI222XL U16877 ( .A0(n20598), .A1(n20537), .B0(n20598), .B1(n20536), .C0(
        n20537), .C1(n20535), .Y(n20595) );
  NOR4BXL U16878 ( .AN(n20534), .B(n20597), .C(n20533), .D(n20532), .Y(n20535)
         );
  INVXL U16879 ( .A(n26172), .Y(n26207) );
  AOI32XL U16880 ( .A0(n24875), .A1(n24874), .A2(n24873), .B0(pool[104]), .B1(
        n24874), .Y(n24901) );
  NOR4XL U16881 ( .A(n24893), .B(n24898), .C(n24890), .D(n24897), .Y(n24875)
         );
  AOI222XL U16882 ( .A0(n24854), .A1(n34999), .B0(n24854), .B1(n35000), .C0(
        n34999), .C1(n35000), .Y(n24874) );
  AOI22XL U16883 ( .A0(n34963), .A1(n35232), .B0(n16663), .B1(n35233), .Y(
        n28286) );
  AOI2BB2XL U16884 ( .B0(n26163), .B1(n26374), .A0N(n26374), .A1N(n26166), .Y(
        n35175) );
  AOI2BB1XL U16885 ( .A0N(pool[134]), .A1N(n35166), .B0(n35165), .Y(n35226) );
  NOR4XL U16886 ( .A(n35125), .B(n35213), .C(n35211), .D(n35124), .Y(n35166)
         );
  NOR2X1 U16887 ( .A(n23261), .B(n23260), .Y(n24458) );
  AOI2BB1XL U16888 ( .A0N(conv_3[504]), .A1N(n32076), .B0(n33918), .Y(n32345)
         );
  NOR2X1 U16889 ( .A(n23517), .B(n23516), .Y(n23772) );
  NAND2X1 U16890 ( .A(n23274), .B(n28467), .Y(n23053) );
  INVX2 U16891 ( .A(n34444), .Y(n27644) );
  NAND2XL U16892 ( .A(n18769), .B(n18768), .Y(n23240) );
  NAND4XL U16893 ( .A(n19092), .B(n19091), .C(n19090), .D(n19089), .Y(n23275)
         );
  AOI222XL U16894 ( .A0(n31392), .A1(n31391), .B0(n31392), .B1(conv_3[349]), 
        .C0(n31391), .C1(conv_3[349]), .Y(n31393) );
  INVXL U16895 ( .A(n34762), .Y(n26717) );
  AOI22X2 U16896 ( .A0(N18471), .A1(n19107), .B0(n22422), .B1(n28467), .Y(
        n19108) );
  INVX2 U16897 ( .A(n34455), .Y(n31871) );
  AOI22XL U16898 ( .A0(n22362), .A1(n23244), .B0(n21100), .B1(n19052), .Y(
        n18949) );
  AOI22XL U16899 ( .A0(n22369), .A1(n23242), .B0(n22370), .B1(n23239), .Y(
        n18948) );
  INVX2 U16900 ( .A(n33535), .Y(n24021) );
  AOI22XL U16901 ( .A0(n22369), .A1(n22169), .B0(n21100), .B1(n23241), .Y(
        n18944) );
  AOI22XL U16902 ( .A0(n22362), .A1(n22172), .B0(n22370), .B1(n23243), .Y(
        n18945) );
  NAND2XL U16903 ( .A(n18745), .B(n18744), .Y(n22122) );
  INVX2 U16904 ( .A(n34740), .Y(n34426) );
  AOI22XL U16905 ( .A0(n23272), .A1(n22152), .B0(n23274), .B1(n22448), .Y(
        n19121) );
  AOI211X2 U16906 ( .A0(n26470), .A1(n22305), .B0(n18968), .C0(n18967), .Y(
        n31418) );
  INVXL U16907 ( .A(n26409), .Y(n34954) );
  INVXL U16908 ( .A(n23053), .Y(n34906) );
  AND2XL U16909 ( .A(n29432), .B(n29431), .Y(n30197) );
  NOR2X1 U16910 ( .A(n29432), .B(n29431), .Y(n30196) );
  NAND2XL U16911 ( .A(n21102), .B(n21101), .Y(n22849) );
  AOI22XL U16912 ( .A0(n22370), .A1(n22202), .B0(n21100), .B1(n22204), .Y(
        n21102) );
  NAND2X1 U16913 ( .A(n19247), .B(n20600), .Y(n18156) );
  NOR2X1 U16914 ( .A(n24945), .B(n24947), .Y(n24943) );
  NOR2X1 U16915 ( .A(n19204), .B(n19205), .Y(n30543) );
  OAI2BB2XL U16916 ( .B0(n22892), .B1(n34989), .A0N(n23092), .A1N(n16755), .Y(
        n22213) );
  NAND2XL U16917 ( .A(n27632), .B(n34019), .Y(n30267) );
  AOI2BB1XL U16918 ( .A0N(conv_1[490]), .A1N(n29992), .B0(n35534), .Y(n30324)
         );
  NAND2XL U16919 ( .A(n27632), .B(n33530), .Y(n35534) );
  NAND2XL U16920 ( .A(n27632), .B(n34706), .Y(n32988) );
  INVXL U16921 ( .A(n34044), .Y(n23394) );
  AOI2BB1XL U16922 ( .A0N(conv_1[53]), .A1N(n27316), .B0(n35309), .Y(n35307)
         );
  AOI2BB1XL U16923 ( .A0N(conv_1[52]), .A1N(n26820), .B0(n35309), .Y(n27316)
         );
  NAND2XL U16924 ( .A(n28739), .B(n34019), .Y(n28706) );
  AOI2BB1XL U16925 ( .A0N(conv_2[489]), .A1N(n27753), .B0(n34130), .Y(n29578)
         );
  AOI2BB1XL U16926 ( .A0N(conv_2[188]), .A1N(n35912), .B0(n30946), .Y(n28657)
         );
  AOI2BB1XL U16927 ( .A0N(conv_2[187]), .A1N(n29885), .B0(n30946), .Y(n35912)
         );
  NAND2XL U16928 ( .A(n34706), .B(n28739), .Y(n30946) );
  NAND2XL U16929 ( .A(n28739), .B(n33990), .Y(n35862) );
  AOI2BB1XL U16930 ( .A0N(conv_3[531]), .A1N(n26369), .B0(n28959), .Y(n27569)
         );
  AOI211XL U16931 ( .A0(n21100), .A1(n34986), .B0(n22245), .C0(n22244), .Y(
        n25688) );
  NAND2XL U16932 ( .A(n32557), .B(n32559), .Y(n32556) );
  AOI2BB1XL U16933 ( .A0N(conv_3[338]), .A1N(n31962), .B0(n31967), .Y(n27590)
         );
  INVXL U16934 ( .A(n31980), .Y(n31967) );
  AOI2BB1XL U16935 ( .A0N(conv_3[190]), .A1N(n31607), .B0(n32207), .Y(n31621)
         );
  AOI21XL U16936 ( .A0(n31602), .A1(conv_3[190]), .B0(n32649), .Y(n31620) );
  NOR2X1 U16937 ( .A(n31609), .B(n31608), .Y(n31602) );
  AOI22XL U16938 ( .A0(n25306), .A1(conv_1[110]), .B0(n16673), .B1(conv_1[140]), .Y(n20015) );
  AOI22XL U16939 ( .A0(n25306), .A1(conv_1[296]), .B0(n22759), .B1(conv_1[281]), .Y(n19960) );
  AOI22XL U16940 ( .A0(n25289), .A1(conv_1[311]), .B0(n22615), .B1(conv_1[326]), .Y(n19959) );
  AOI22XL U16941 ( .A0(n36246), .A1(n22596), .B0(n22595), .B1(n22765), .Y(
        n28534) );
  AOI22XL U16942 ( .A0(n25299), .A1(conv_2[157]), .B0(n22615), .B1(conv_2[202]), .Y(n20932) );
  AOI22XL U16943 ( .A0(n22762), .A1(conv_2[352]), .B0(n22615), .B1(conv_2[382]), .Y(n20947) );
  AOI22XL U16944 ( .A0(n25299), .A1(conv_2[277]), .B0(n22615), .B1(conv_2[322]), .Y(n20937) );
  AOI22XL U16945 ( .A0(n36246), .A1(n26009), .B0(n26027), .B1(n22743), .Y(
        n26015) );
  NOR2X1 U16946 ( .A(n19284), .B(n19283), .Y(n21245) );
  AOI22XL U16947 ( .A0(n22759), .A1(conv_3[36]), .B0(n22615), .B1(conv_3[81]), 
        .Y(n19324) );
  AOI22XL U16948 ( .A0(n34963), .A1(n21362), .B0(conv_3[220]), .B1(n16744), 
        .Y(n20482) );
  AOI22XL U16949 ( .A0(n16666), .A1(conv_3[56]), .B0(n25289), .B1(conv_3[71]), 
        .Y(n19295) );
  AOI22XL U16950 ( .A0(n22759), .A1(conv_3[41]), .B0(n22615), .B1(conv_3[86]), 
        .Y(n19296) );
  AOI22XL U16951 ( .A0(n22759), .A1(conv_3[101]), .B0(n22615), .B1(conv_3[146]), .Y(n19298) );
  AOI22XL U16952 ( .A0(n25289), .A1(conv_1[371]), .B0(n22759), .B1(conv_1[341]), .Y(n19962) );
  AOI22XL U16953 ( .A0(n25306), .A1(conv_1[356]), .B0(n22615), .B1(conv_1[386]), .Y(n19961) );
  AOI22XL U16954 ( .A0(n25306), .A1(conv_1[116]), .B0(n22615), .B1(conv_1[146]), .Y(n19956) );
  AOI211XL U16955 ( .A0(conv_1[175]), .A1(n25306), .B0(n19922), .C0(n19921), 
        .Y(n21654) );
  AOI22XL U16956 ( .A0(n25306), .A1(conv_1[56]), .B0(n22759), .B1(conv_1[41]), 
        .Y(n19957) );
  AOI22XL U16957 ( .A0(n16662), .A1(conv_1[71]), .B0(n22615), .B1(conv_1[86]), 
        .Y(n19958) );
  AOI22XL U16958 ( .A0(n36246), .A1(n22595), .B0(n22596), .B1(n22743), .Y(
        n21677) );
  AOI22XL U16959 ( .A0(n25306), .A1(conv_1[176]), .B0(n16662), .B1(conv_1[191]), .Y(n19952) );
  AOI22XL U16960 ( .A0(n22759), .A1(conv_1[161]), .B0(n22615), .B1(conv_1[206]), .Y(n19953) );
  AOI22XL U16961 ( .A0(n34992), .A1(n21674), .B0(n34963), .B1(n21687), .Y(
        n19966) );
  AOI22XL U16962 ( .A0(n34963), .A1(n28515), .B0(n26262), .B1(n28513), .Y(
        n25352) );
  AOI22XL U16963 ( .A0(n25306), .A1(conv_1[321]), .B0(n25299), .B1(conv_1[306]), .Y(n22470) );
  AOI22XL U16964 ( .A0(n25306), .A1(conv_1[22]), .B0(n16673), .B1(conv_1[52]), 
        .Y(n22624) );
  AOI22XL U16965 ( .A0(n36246), .A1(n22627), .B0(n22626), .B1(n22743), .Y(
        n28470) );
  AOI211XL U16966 ( .A0(conv_1[215]), .A1(n25289), .B0(n22573), .C0(n22572), 
        .Y(n28489) );
  AOI22XL U16967 ( .A0(n25306), .A1(conv_1[80]), .B0(n16673), .B1(conv_1[110]), 
        .Y(n22576) );
  AOI22XL U16968 ( .A0(n25306), .A1(conv_1[141]), .B0(n16662), .B1(conv_1[156]), .Y(n22468) );
  AOI22XL U16969 ( .A0(n25306), .A1(conv_1[142]), .B0(n25299), .B1(conv_1[127]), .Y(n22609) );
  AOI22XL U16970 ( .A0(n25306), .A1(conv_1[82]), .B0(n16662), .B1(conv_1[97]), 
        .Y(n22618) );
  AOI22XL U16971 ( .A0(n25306), .A1(conv_1[382]), .B0(n16662), .B1(conv_1[397]), .Y(n22619) );
  AOI211XL U16972 ( .A0(conv_1[232]), .A1(n22615), .B0(n22614), .C0(n22613), 
        .Y(n28472) );
  AOI211XL U16973 ( .A0(n22759), .A1(conv_1[6]), .B0(n22462), .C0(n22461), .Y(
        n28503) );
  AOI22XL U16974 ( .A0(n36246), .A1(n22464), .B0(n22463), .B1(n21358), .Y(
        n28511) );
  AND2XL U16975 ( .A(n22543), .B(n22542), .Y(n28440) );
  AOI22XL U16976 ( .A0(n25306), .A1(conv_1[143]), .B0(n22690), .B1(conv_1[128]), .Y(n22542) );
  AOI211XL U16977 ( .A0(conv_2[174]), .A1(n25306), .B0(n20874), .C0(n20873), 
        .Y(n25999) );
  AOI22XL U16978 ( .A0(n16662), .A1(conv_2[71]), .B0(n22615), .B1(conv_2[86]), 
        .Y(n20888) );
  OAI211XL U16979 ( .A0(n36246), .A1(n25960), .B0(n28528), .C0(n25959), .Y(
        n25961) );
  NAND2XL U16980 ( .A(n36246), .B(n25958), .Y(n25959) );
  OAI211XL U16981 ( .A0(n36246), .A1(n26011), .B0(n28528), .C0(n26010), .Y(
        n26012) );
  NAND2XL U16982 ( .A(n36246), .B(n26009), .Y(n26010) );
  AOI211XL U16983 ( .A0(conv_2[131]), .A1(n25289), .B0(n20896), .C0(n20895), 
        .Y(n26014) );
  AOI22XL U16984 ( .A0(n22762), .A1(conv_2[176]), .B0(n22615), .B1(conv_2[206]), .Y(n20897) );
  AOI22XL U16985 ( .A0(n25306), .A1(conv_2[58]), .B0(n22759), .B1(conv_2[43]), 
        .Y(n21064) );
  AOI22XL U16986 ( .A0(n16662), .A1(conv_2[73]), .B0(n22615), .B1(conv_2[88]), 
        .Y(n21065) );
  AOI22XL U16987 ( .A0(n21011), .A1(conv_2[354]), .B0(n22615), .B1(conv_2[384]), .Y(n20869) );
  AOI211XL U16988 ( .A0(conv_2[129]), .A1(n25289), .B0(n20864), .C0(n20863), 
        .Y(n25998) );
  NOR2X1 U16989 ( .A(n22717), .B(n30944), .Y(n20864) );
  AOI22XL U16990 ( .A0(n25289), .A1(conv_2[396]), .B0(n22690), .B1(conv_2[366]), .Y(n18281) );
  AOI22XL U16991 ( .A0(n25289), .A1(conv_2[336]), .B0(n16673), .B1(conv_2[351]), .Y(n18283) );
  AOI211XL U16992 ( .A0(n16673), .A1(conv_2[232]), .B0(n18306), .C0(n18305), 
        .Y(n25148) );
  AOI22XL U16993 ( .A0(n25289), .A1(conv_2[96]), .B0(n25299), .B1(conv_2[66]), 
        .Y(n18290) );
  AOI22XL U16994 ( .A0(n25289), .A1(conv_2[156]), .B0(n22759), .B1(conv_2[126]), .Y(n18285) );
  AOI22XL U16995 ( .A0(n36246), .A1(n25915), .B0(n20946), .B1(n21358), .Y(
        n25147) );
  AOI22XL U16996 ( .A0(n25289), .A1(conv_2[37]), .B0(n16673), .B1(conv_2[52]), 
        .Y(n18302) );
  AOI22XL U16997 ( .A0(n36246), .A1(n21879), .B0(n21880), .B1(n21688), .Y(
        n25519) );
  AOI211XL U16998 ( .A0(conv_2[65]), .A1(n22616), .B0(n18242), .C0(n18241), 
        .Y(n25514) );
  AOI211XL U16999 ( .A0(n25289), .A1(conv_2[155]), .B0(n18236), .C0(n18235), 
        .Y(n25513) );
  NOR2X1 U17000 ( .A(n24039), .B(n29838), .Y(n18236) );
  AOI22XL U17001 ( .A0(n36246), .A1(n25955), .B0(n25958), .B1(n22713), .Y(
        n25542) );
  AOI22XL U17002 ( .A0(n25289), .A1(conv_2[97]), .B0(n16673), .B1(conv_2[112]), 
        .Y(n18303) );
  AOI22XL U17003 ( .A0(n25289), .A1(conv_2[101]), .B0(n25299), .B1(conv_2[71]), 
        .Y(n18335) );
  NOR2X1 U17004 ( .A(n18750), .B(n31459), .Y(n19286) );
  AOI22XL U17005 ( .A0(n16662), .A1(conv_3[311]), .B0(n22615), .B1(conv_3[326]), .Y(n19294) );
  AOI22XL U17006 ( .A0(n36246), .A1(n20473), .B0(n21313), .B1(n22743), .Y(
        n21305) );
  AOI22XL U17007 ( .A0(n22759), .A1(conv_3[158]), .B0(n22615), .B1(conv_3[203]), .Y(n19406) );
  AOI22XL U17008 ( .A0(n22759), .A1(conv_3[98]), .B0(n22615), .B1(conv_3[143]), 
        .Y(n19408) );
  AOI22XL U17009 ( .A0(n16666), .A1(conv_3[353]), .B0(n22615), .B1(conv_3[383]), .Y(n19411) );
  AOI22XL U17010 ( .A0(n28528), .A1(n35052), .B0(n34963), .B1(n26193), .Y(
        n26194) );
  AOI22XL U17011 ( .A0(n36246), .A1(n21226), .B0(n21213), .B1(n22713), .Y(
        n35090) );
  AOI22XL U17012 ( .A0(n36246), .A1(n21263), .B0(n21269), .B1(n22713), .Y(
        n35070) );
  NOR2X1 U17013 ( .A(n22612), .B(n31249), .Y(n18552) );
  AOI22XL U17014 ( .A0(n20978), .A1(conv_3[142]), .B0(n22615), .B1(conv_3[172]), .Y(n18537) );
  AOI22XL U17015 ( .A0(n16662), .A1(conv_3[217]), .B0(n22615), .B1(conv_3[232]), .Y(n18530) );
  AOI22XL U17016 ( .A0(n16666), .A1(conv_3[382]), .B0(n22615), .B1(conv_3[412]), .Y(n18528) );
  AOI22XL U17017 ( .A0(n36246), .A1(n21313), .B0(n20473), .B1(n22713), .Y(
        n35114) );
  NOR4XL U17018 ( .A(n17835), .B(n17834), .C(n17833), .D(n17832), .Y(n17911)
         );
  NOR4XL U17019 ( .A(n17908), .B(n17907), .C(n17906), .D(n17905), .Y(n17909)
         );
  NOR4XL U17020 ( .A(n17862), .B(n17861), .C(n17860), .D(n17859), .Y(n17910)
         );
  NOR2X1 U17021 ( .A(n20755), .B(n18109), .Y(n17801) );
  NOR3XL U17022 ( .A(n18103), .B(n18102), .C(n18101), .Y(n18104) );
  NOR3XL U17023 ( .A(n17959), .B(n17958), .C(n17957), .Y(n17960) );
  AOI221XL U17024 ( .A0(n19611), .A1(n19614), .B0(n18037), .B1(n19613), .C0(
        n19612), .Y(n18070) );
  INVXL U17025 ( .A(n19612), .Y(n19622) );
  INVXL U17026 ( .A(n18070), .Y(n19616) );
  INVXL U17027 ( .A(n17989), .Y(n19689) );
  AOI22XL U17028 ( .A0(n25306), .A1(conv_1[166]), .B0(n16673), .B1(conv_1[196]), .Y(n19841) );
  AOI22XL U17029 ( .A0(n16662), .A1(conv_2[61]), .B0(n22615), .B1(conv_2[76]), 
        .Y(n21016) );
  AOI22XL U17030 ( .A0(n25299), .A1(conv_2[271]), .B0(n22615), .B1(conv_2[316]), .Y(n21006) );
  NAND2XL U17031 ( .A(n21013), .B(n21012), .Y(n25882) );
  AOI22XL U17032 ( .A0(n21011), .A1(conv_2[346]), .B0(n22615), .B1(conv_2[376]), .Y(n21013) );
  NAND2XL U17033 ( .A(n19509), .B(n19508), .Y(n21158) );
  AOI22XL U17034 ( .A0(n22690), .A1(conv_3[31]), .B0(n22615), .B1(conv_3[76]), 
        .Y(n19508) );
  AOI22XL U17035 ( .A0(n16662), .A1(conv_3[181]), .B0(n22615), .B1(conv_3[196]), .Y(n19504) );
  AOI22XL U17036 ( .A0(n16666), .A1(conv_3[286]), .B0(n22615), .B1(conv_3[316]), .Y(n19510) );
  AOI22XL U17037 ( .A0(n16666), .A1(conv_3[346]), .B0(n22615), .B1(conv_3[376]), .Y(n19507) );
  AOI22XL U17038 ( .A0(n25289), .A1(conv_3[121]), .B0(n22615), .B1(conv_3[136]), .Y(n19503) );
  AOI22XL U17039 ( .A0(n25306), .A1(conv_1[167]), .B0(n16662), .B1(conv_1[182]), .Y(n19822) );
  AOI22XL U17040 ( .A0(n25306), .A1(conv_2[287]), .B0(n22615), .B1(conv_2[317]), .Y(n20991) );
  AOI22XL U17041 ( .A0(n25299), .A1(conv_2[92]), .B0(n22615), .B1(conv_2[137]), 
        .Y(n20986) );
  AOI22XL U17042 ( .A0(n25306), .A1(conv_2[107]), .B0(n25289), .B1(conv_2[122]), .Y(n20987) );
  AOI22XL U17043 ( .A0(n16662), .A1(conv_2[62]), .B0(n22615), .B1(conv_2[77]), 
        .Y(n20989) );
  AOI22XL U17044 ( .A0(n25306), .A1(conv_2[347]), .B0(n22615), .B1(conv_2[377]), .Y(n20984) );
  AOI22XL U17045 ( .A0(n19007), .A1(filter_2[25]), .B0(n16676), .B1(
        filter_2[37]), .Y(n18910) );
  AOI22XL U17046 ( .A0(n36246), .A1(n22644), .B0(n22643), .B1(n22743), .Y(
        n25373) );
  INVXL U17047 ( .A(n25373), .Y(n26384) );
  AOI22XL U17048 ( .A0(n19006), .A1(filter_1[8]), .B0(n19007), .B1(
        filter_1[26]), .Y(n18832) );
  AOI22XL U17049 ( .A0(n19004), .A1(filter_1[32]), .B0(n16676), .B1(
        filter_1[38]), .Y(n18831) );
  AND2XL U17050 ( .A(n22391), .B(n26698), .Y(n22392) );
  AOI22XL U17051 ( .A0(n25306), .A1(conv_2[348]), .B0(n22615), .B1(conv_2[378]), .Y(n20966) );
  AOI22XL U17052 ( .A0(n25306), .A1(conv_2[168]), .B0(n25289), .B1(conv_2[183]), .Y(n20962) );
  AOI22XL U17053 ( .A0(n25299), .A1(conv_2[153]), .B0(n22615), .B1(conv_2[198]), .Y(n20963) );
  AOI22XL U17054 ( .A0(n36246), .A1(n21818), .B0(n25836), .B1(n22765), .Y(
        n24956) );
  AOI22XL U17055 ( .A0(n25289), .A1(conv_3[63]), .B0(n18240), .B1(conv_3[78]), 
        .Y(n19457) );
  AOI22XL U17056 ( .A0(n25289), .A1(conv_3[303]), .B0(n18240), .B1(conv_3[318]), .Y(n19462) );
  AOI22XL U17057 ( .A0(n25289), .A1(conv_3[363]), .B0(n22615), .B1(conv_3[378]), .Y(n19459) );
  AOI22XL U17058 ( .A0(n19009), .A1(filter_3[20]), .B0(n19007), .B1(
        filter_3[26]), .Y(n18992) );
  AOI22XL U17059 ( .A0(n19006), .A1(filter_3[8]), .B0(n19004), .B1(
        filter_3[32]), .Y(n18993) );
  OAI222XL U17060 ( .A0(n30771), .A1(n22612), .B0(n36246), .B1(n22498), .C0(
        n30778), .C1(n24039), .Y(n26413) );
  AOI22XL U17061 ( .A0(n25306), .A1(conv_1[319]), .B0(n22616), .B1(conv_1[304]), .Y(n22502) );
  AOI22XL U17062 ( .A0(n25306), .A1(conv_1[379]), .B0(n16673), .B1(conv_1[409]), .Y(n22504) );
  AOI22XL U17063 ( .A0(n16662), .A1(conv_2[124]), .B0(n22615), .B1(conv_2[139]), .Y(n20773) );
  AOI22XL U17064 ( .A0(n25299), .A1(conv_2[274]), .B0(n22615), .B1(conv_2[319]), .Y(n20780) );
  AOI22XL U17065 ( .A0(n16662), .A1(conv_2[64]), .B0(n22615), .B1(conv_2[79]), 
        .Y(n20777) );
  AOI22XL U17066 ( .A0(n22762), .A1(conv_2[349]), .B0(n22615), .B1(conv_2[379]), .Y(n20775) );
  AOI22XL U17067 ( .A0(n25289), .A1(conv_2[154]), .B0(n16673), .B1(conv_2[169]), .Y(n18252) );
  AOI222X1 U17068 ( .A0(n29002), .A1(conv_2[168]), .B0(n29002), .B1(n29001), 
        .C0(conv_2[168]), .C1(n29001), .Y(n29003) );
  AOI22XL U17069 ( .A0(n16662), .A1(conv_3[184]), .B0(n22615), .B1(conv_3[199]), .Y(n19371) );
  NOR2X1 U17070 ( .A(n36244), .B(n24828), .Y(n18498) );
  AOI22XL U17071 ( .A0(n18658), .A1(conv_3[364]), .B0(n22615), .B1(conv_3[409]), .Y(n18501) );
  AOI22XL U17072 ( .A0(n34963), .A1(n28526), .B0(n26276), .B1(n28527), .Y(
        n25367) );
  AOI22XL U17073 ( .A0(n36246), .A1(n22721), .B0(n22720), .B1(n21358), .Y(
        n28421) );
  AOI22XL U17074 ( .A0(n25306), .A1(conv_1[389]), .B0(n25299), .B1(conv_1[374]), .Y(n22708) );
  AOI2BB1XL U17075 ( .A0N(conv_1[124]), .A1N(n30753), .B0(n30754), .Y(n23650)
         );
  INVX2 U17076 ( .A(n16725), .Y(n16715) );
  AOI22XL U17077 ( .A0(n25306), .A1(conv_2[358]), .B0(n18240), .B1(conv_2[388]), .Y(n21062) );
  NAND2XL U17078 ( .A(n36246), .B(n22012), .Y(n26089) );
  NAND2XL U17079 ( .A(n36246), .B(n21976), .Y(n25815) );
  AOI211XL U17080 ( .A0(conv_2[299]), .A1(n25306), .B0(n20761), .C0(n20760), 
        .Y(n25814) );
  AOI22XL U17081 ( .A0(n28528), .A1(n25648), .B0(n34963), .B1(n25657), .Y(
        n24113) );
  AOI22XL U17082 ( .A0(n25306), .A1(conv_2[375]), .B0(n16662), .B1(conv_2[390]), .Y(n24031) );
  AOI2BB1XL U17083 ( .A0N(conv_2[319]), .A1N(n28864), .B0(n28865), .Y(n23106)
         );
  AOI2BB1XL U17084 ( .A0N(conv_2[214]), .A1N(n28876), .B0(n28877), .Y(n28665)
         );
  NOR2X1 U17085 ( .A(n29166), .B(n26085), .Y(n19448) );
  AOI22XL U17086 ( .A0(n16666), .A1(conv_3[57]), .B0(n25289), .B1(conv_3[72]), 
        .Y(n19549) );
  AOI211XL U17087 ( .A0(n34963), .A1(n35040), .B0(n24870), .C0(n24869), .Y(
        n24871) );
  AOI22XL U17088 ( .A0(n36246), .A1(n21388), .B0(n20538), .B1(n22743), .Y(
        n35169) );
  NOR2XL U17089 ( .A(n31691), .B(n27764), .Y(n23261) );
  NAND2XL U17090 ( .A(n18743), .B(n18742), .Y(n19050) );
  NAND2XL U17091 ( .A(n18733), .B(n18732), .Y(n22169) );
  NOR2X1 U17092 ( .A(n30195), .B(n31691), .Y(n29432) );
  AOI22XL U17093 ( .A0(n19006), .A1(filter_3[10]), .B0(n19007), .B1(
        filter_3[28]), .Y(n18982) );
  AOI2BB1XL U17094 ( .A0N(n20618), .A1N(n33563), .B0(n20617), .Y(n33075) );
  OAI2BB1XL U17095 ( .A0N(weight_2[48]), .A1N(n18049), .B0(n18009), .Y(n18010)
         );
  OAI221X1 U17096 ( .A0(n18054), .A1(n24561), .B0(n18053), .B1(n24560), .C0(
        n28398), .Y(n28397) );
  OAI221X1 U17097 ( .A0(n17984), .A1(n24544), .B0(n17983), .B1(n24543), .C0(
        n28211), .Y(n28210) );
  NAND2X1 U17098 ( .A(n19243), .B(ns[0]), .Y(n19610) );
  AOI22XL U17099 ( .A0(n25306), .A1(conv_1[106]), .B0(n16673), .B1(conv_1[136]), .Y(n19838) );
  NAND2XL U17100 ( .A(n19846), .B(n19845), .Y(n21505) );
  AOI22XL U17101 ( .A0(n25306), .A1(conv_1[346]), .B0(n16673), .B1(conv_1[376]), .Y(n19845) );
  AOI22XL U17102 ( .A0(n25289), .A1(conv_1[361]), .B0(n22690), .B1(conv_1[331]), .Y(n19846) );
  AOI22XL U17103 ( .A0(n36246), .A1(n22682), .B0(n22683), .B1(n22713), .Y(
        n21501) );
  AOI22XL U17104 ( .A0(n25306), .A1(conv_1[286]), .B0(n16662), .B1(conv_1[301]), .Y(n19844) );
  AOI211XL U17105 ( .A0(conv_1[61]), .A1(n25289), .B0(n19840), .C0(n19839), 
        .Y(n21497) );
  AOI22XL U17106 ( .A0(n36246), .A1(n22683), .B0(n22682), .B1(n22765), .Y(
        n25400) );
  AND2XL U17107 ( .A(n22692), .B(n22691), .Y(n25396) );
  AOI22XL U17108 ( .A0(n16716), .A1(conv_1[331]), .B0(n22690), .B1(conv_1[301]), .Y(n22691) );
  NAND2XL U17109 ( .A(n33873), .B(n27429), .Y(n22292) );
  NAND2XL U17110 ( .A(n21003), .B(n21002), .Y(n25880) );
  AOI22XL U17111 ( .A0(n16662), .A1(conv_2[121]), .B0(n22615), .B1(conv_2[136]), .Y(n21003) );
  NAND2XL U17112 ( .A(n36246), .B(n34963), .Y(n21004) );
  NAND2XL U17113 ( .A(n21015), .B(n21014), .Y(n25870) );
  AOI22XL U17114 ( .A0(n22762), .A1(conv_2[166]), .B0(n22690), .B1(conv_2[151]), .Y(n21014) );
  AOI22XL U17115 ( .A0(n34963), .A1(n25877), .B0(n24056), .B1(n25878), .Y(
        n21851) );
  AOI22XL U17116 ( .A0(n25289), .A1(conv_2[31]), .B0(n16673), .B1(conv_2[46]), 
        .Y(n18382) );
  AOI22XL U17117 ( .A0(n25289), .A1(conv_2[151]), .B0(n22690), .B1(conv_2[121]), .Y(n18390) );
  AOI22XL U17118 ( .A0(n25289), .A1(conv_2[211]), .B0(n16673), .B1(conv_2[226]), .Y(n18392) );
  INVXL U17119 ( .A(n24709), .Y(n25113) );
  AOI22XL U17120 ( .A0(n36246), .A1(n25874), .B0(n21849), .B1(n21688), .Y(
        n24971) );
  OAI222XL U17121 ( .A0(n24554), .A1(n22612), .B0(n36246), .B1(n25873), .C0(
        n30305), .C1(n18750), .Y(n25487) );
  AOI22XL U17122 ( .A0(n25306), .A1(conv_2[376]), .B0(n16662), .B1(conv_2[391]), .Y(n18386) );
  AOI22XL U17123 ( .A0(n36246), .A1(n21148), .B0(n21147), .B1(n22713), .Y(
        n21155) );
  AOI22XL U17124 ( .A0(n16667), .A1(n21154), .B0(n34963), .B1(n21158), .Y(
        n20446) );
  AOI22XL U17125 ( .A0(n36246), .A1(n21147), .B0(n21148), .B1(n21688), .Y(
        n35153) );
  INVXL U17126 ( .A(n31376), .Y(n19015) );
  AOI22XL U17127 ( .A0(n25306), .A1(conv_1[347]), .B0(n22690), .B1(conv_1[332]), .Y(n19814) );
  AOI22XL U17128 ( .A0(n25306), .A1(conv_1[287]), .B0(n16662), .B1(conv_1[302]), .Y(n19818) );
  AOI22XL U17129 ( .A0(n25306), .A1(conv_1[47]), .B0(n22759), .B1(conv_1[32]), 
        .Y(n19815) );
  AOI22XL U17130 ( .A0(n25306), .A1(conv_1[107]), .B0(n22690), .B1(conv_1[92]), 
        .Y(n19819) );
  AOI22XL U17131 ( .A0(n34963), .A1(n21516), .B0(n34961), .B1(n21521), .Y(
        n19824) );
  NOR2X1 U17132 ( .A(n26556), .B(n25123), .Y(n22667) );
  AOI211XL U17133 ( .A0(n25399), .A1(n25387), .B0(n25386), .C0(n25385), .Y(
        n28428) );
  AOI22XL U17134 ( .A0(n36245), .A1(n25387), .B0(n25384), .B1(n26374), .Y(
        n26557) );
  INVXL U17135 ( .A(n24618), .Y(n26562) );
  AOI22XL U17136 ( .A0(n36246), .A1(n22657), .B0(n22656), .B1(n22765), .Y(
        n24618) );
  AND2XL U17137 ( .A(n22671), .B(n22670), .Y(n26555) );
  NOR2X1 U17138 ( .A(n36244), .B(n24618), .Y(n22673) );
  NOR2X1 U17139 ( .A(n33399), .B(n33398), .Y(n33400) );
  NOR2X1 U17140 ( .A(n34521), .B(n22940), .Y(n22941) );
  AOI22XL U17141 ( .A0(n34963), .A1(n25858), .B0(n35234), .B1(n25856), .Y(
        n21835) );
  AOI22XL U17142 ( .A0(n25299), .A1(conv_2[152]), .B0(n22615), .B1(conv_2[197]), .Y(n20980) );
  AOI22XL U17143 ( .A0(n25306), .A1(conv_2[17]), .B0(n16662), .B1(conv_2[32]), 
        .Y(n18371) );
  AND2XL U17144 ( .A(n18370), .B(n18369), .Y(n25124) );
  AOI22XL U17145 ( .A0(n25289), .A1(conv_2[92]), .B0(n22690), .B1(conv_2[62]), 
        .Y(n18370) );
  AOI22XL U17146 ( .A0(n36246), .A1(n20981), .B0(n25854), .B1(n22743), .Y(
        n25119) );
  AOI22XL U17147 ( .A0(n25306), .A1(conv_2[197]), .B0(n16662), .B1(conv_2[212]), .Y(n18368) );
  AOI22XL U17148 ( .A0(n25289), .A1(conv_2[152]), .B0(n16673), .B1(conv_2[167]), .Y(n18366) );
  AOI22XL U17149 ( .A0(n25306), .A1(conv_2[317]), .B0(n22690), .B1(conv_2[302]), .Y(n18377) );
  NAND2XL U17150 ( .A(n23348), .B(n31090), .Y(n23350) );
  NAND2XL U17151 ( .A(n23475), .B(n23946), .Y(n23477) );
  AOI22XL U17152 ( .A0(n22690), .A1(conv_3[332]), .B0(n22615), .B1(conv_3[377]), .Y(n19483) );
  AOI211XL U17153 ( .A0(conv_3[392]), .A1(n21749), .B0(n21183), .C0(n21182), 
        .Y(n21184) );
  AOI22XL U17154 ( .A0(n22690), .A1(conv_3[272]), .B0(n22615), .B1(conv_3[317]), .Y(n19493) );
  AOI22XL U17155 ( .A0(n25289), .A1(conv_3[62]), .B0(n22690), .B1(conv_3[32]), 
        .Y(n19472) );
  AOI22XL U17156 ( .A0(n16666), .A1(conv_3[47]), .B0(n22615), .B1(conv_3[77]), 
        .Y(n19473) );
  AOI22XL U17157 ( .A0(n22690), .A1(conv_3[92]), .B0(n22615), .B1(conv_3[137]), 
        .Y(n19484) );
  AOI22XL U17158 ( .A0(n36246), .A1(n19470), .B0(n20432), .B1(n22713), .Y(
        n28278) );
  AOI22XL U17159 ( .A0(n25289), .A1(conv_3[152]), .B0(n16673), .B1(conv_3[167]), .Y(n18622) );
  AOI22XL U17160 ( .A0(n22762), .A1(conv_3[317]), .B0(n22615), .B1(conv_3[347]), .Y(n18617) );
  AOI22XL U17161 ( .A0(n22762), .A1(conv_3[377]), .B0(n22615), .B1(conv_3[407]), .Y(n18615) );
  NAND2XL U17162 ( .A(n36246), .B(n22643), .Y(n20206) );
  AOI22XL U17163 ( .A0(n34963), .A1(n21480), .B0(n34961), .B1(n21484), .Y(
        n19802) );
  OR2XL U17164 ( .A(n17173), .B(n23053), .Y(n22008) );
  NOR2X1 U17165 ( .A(n25373), .B(n16721), .Y(n26382) );
  AOI22XL U17166 ( .A0(n16755), .A1(n26382), .B0(n34963), .B1(n26537), .Y(
        n26383) );
  INVXL U17167 ( .A(n25375), .Y(n24615) );
  NOR2X1 U17168 ( .A(n35498), .B(n23504), .Y(n28966) );
  NOR2X1 U17169 ( .A(n35498), .B(n28721), .Y(n23467) );
  NOR2X1 U17170 ( .A(n35272), .B(n33491), .Y(n22429) );
  NOR2X1 U17171 ( .A(n35498), .B(n34715), .Y(n31370) );
  NOR2X1 U17172 ( .A(n22392), .B(n22393), .Y(n26684) );
  AND2XL U17173 ( .A(n22393), .B(n22392), .Y(n26685) );
  AOI22XL U17174 ( .A0(n25306), .A1(conv_2[288]), .B0(n22615), .B1(conv_2[318]), .Y(n20960) );
  NAND2XL U17175 ( .A(n21004), .B(n21311), .Y(n21753) );
  AOI22XL U17176 ( .A0(n25306), .A1(conv_2[108]), .B0(n16662), .B1(conv_2[123]), .Y(n20965) );
  AOI22XL U17177 ( .A0(n25299), .A1(conv_2[93]), .B0(n22615), .B1(conv_2[138]), 
        .Y(n20964) );
  NAND2XL U17178 ( .A(n36246), .B(n16659), .Y(n25987) );
  AOI22XL U17179 ( .A0(n34963), .A1(n25842), .B0(n34961), .B1(n25841), .Y(
        n21820) );
  AOI22XL U17180 ( .A0(n25306), .A1(conv_2[18]), .B0(n22690), .B1(conv_2[3]), 
        .Y(n18348) );
  AOI22XL U17181 ( .A0(n25306), .A1(conv_2[138]), .B0(n16673), .B1(conv_2[168]), .Y(n18355) );
  AOI22XL U17182 ( .A0(n25306), .A1(conv_2[318]), .B0(n16673), .B1(conv_2[348]), .Y(n18353) );
  AOI2BB1XL U17183 ( .A0N(conv_2[392]), .A1N(n30343), .B0(n30344), .Y(n24448)
         );
  NOR2X1 U17184 ( .A(n34703), .B(n35856), .Y(n28652) );
  NOR2X1 U17185 ( .A(n23112), .B(n23111), .Y(n23267) );
  NOR2X1 U17186 ( .A(n35856), .B(n34715), .Y(n27139) );
  NOR2XL U17187 ( .A(n35856), .B(n31418), .Y(n26742) );
  AOI22XL U17188 ( .A0(n25289), .A1(conv_3[123]), .B0(n22690), .B1(conv_3[93]), 
        .Y(n19454) );
  AOI22XL U17189 ( .A0(n28528), .A1(n21135), .B0(n34963), .B1(n21134), .Y(
        n20423) );
  NAND2XL U17190 ( .A(n34827), .B(n21991), .Y(n21959) );
  AOI22XL U17191 ( .A0(n25306), .A1(conv_3[198]), .B0(n25289), .B1(conv_3[213]), .Y(n18598) );
  AOI211XL U17192 ( .A0(n25399), .A1(n25699), .B0(n18607), .C0(n18606), .Y(
        n26175) );
  AOI22XL U17193 ( .A0(n36246), .A1(n20422), .B0(n21123), .B1(n21688), .Y(
        n26171) );
  AOI211XL U17194 ( .A0(n22370), .A1(n35128), .B0(n35129), .C0(n24849), .Y(
        n28274) );
  NOR2X1 U17195 ( .A(n36245), .B(n24848), .Y(n24849) );
  AOI22XL U17196 ( .A0(n18658), .A1(conv_3[123]), .B0(n22615), .B1(conv_3[168]), .Y(n18600) );
  INVXL U17197 ( .A(n35231), .Y(n35143) );
  AOI222XL U17198 ( .A0(n30780), .A1(conv_3[467]), .B0(n30780), .B1(n30779), 
        .C0(conv_3[467]), .C1(n30779), .Y(n19017) );
  NOR2X1 U17199 ( .A(n29426), .B(n23504), .Y(n23506) );
  NOR2X1 U17200 ( .A(n29426), .B(n33994), .Y(n23492) );
  AOI222XL U17201 ( .A0(n30575), .A1(conv_3[257]), .B0(n30575), .B1(n30574), 
        .C0(conv_3[257]), .C1(n30574), .Y(n22111) );
  AOI222XL U17202 ( .A0(n30824), .A1(conv_3[92]), .B0(n30824), .B1(n30823), 
        .C0(conv_3[92]), .C1(n30823), .Y(n22874) );
  OR2XL U17203 ( .A(n23898), .B(n23897), .Y(n34108) );
  AOI22XL U17204 ( .A0(n25306), .A1(conv_1[19]), .B0(n25299), .B1(conv_1[4]), 
        .Y(n22514) );
  AOI22XL U17205 ( .A0(n25306), .A1(conv_1[199]), .B0(n16662), .B1(conv_1[214]), .Y(n22506) );
  AOI22XL U17206 ( .A0(n36246), .A1(n22510), .B0(n22509), .B1(n22743), .Y(
        n26410) );
  AOI22XL U17207 ( .A0(n25306), .A1(conv_1[139]), .B0(n16662), .B1(conv_1[154]), .Y(n22508) );
  AOI22XL U17208 ( .A0(n25306), .A1(conv_1[79]), .B0(n16662), .B1(conv_1[94]), 
        .Y(n22513) );
  NOR2X1 U17209 ( .A(n35500), .B(n27735), .Y(n27219) );
  INVXL U17210 ( .A(n18852), .Y(n18853) );
  AOI222XL U17211 ( .A0(n26952), .A1(conv_1[468]), .B0(n26952), .B1(n26951), 
        .C0(conv_1[468]), .C1(n26951), .Y(n18852) );
  NOR2X1 U17212 ( .A(n35500), .B(n27860), .Y(n18854) );
  NOR2X1 U17213 ( .A(n35500), .B(n32016), .Y(n27636) );
  AND2XL U17214 ( .A(n24318), .B(n24317), .Y(n30282) );
  NOR2X1 U17215 ( .A(n35500), .B(n24021), .Y(n24439) );
  NOR2X1 U17216 ( .A(n35500), .B(n28660), .Y(n23998) );
  NOR2XL U17217 ( .A(n35500), .B(n22257), .Y(n24496) );
  NOR2X1 U17218 ( .A(n35500), .B(n23296), .Y(n24008) );
  AND2XL U17219 ( .A(n23649), .B(n23648), .Y(n30753) );
  AND2XL U17220 ( .A(n26513), .B(n26512), .Y(n26921) );
  NOR2XL U17221 ( .A(n35500), .B(n31418), .Y(n27405) );
  AOI2BB1XL U17222 ( .A0N(conv_1[18]), .A1N(n27356), .B0(n27357), .Y(n26503)
         );
  NOR2X1 U17223 ( .A(n30195), .B(n35500), .Y(n26504) );
  AOI22XL U17224 ( .A0(n25289), .A1(conv_2[34]), .B0(n16673), .B1(conv_2[49]), 
        .Y(n18253) );
  AOI22XL U17225 ( .A0(n25289), .A1(conv_2[94]), .B0(n22759), .B1(conv_2[64]), 
        .Y(n18247) );
  AOI22XL U17226 ( .A0(n25306), .A1(conv_2[319]), .B0(n16662), .B1(conv_2[334]), .Y(n18259) );
  AOI22XL U17227 ( .A0(n36246), .A1(n25936), .B0(n21866), .B1(n22765), .Y(
        n25501) );
  AOI2BB1XL U17228 ( .A0N(conv_2[438]), .A1N(n29553), .B0(n29554), .Y(n27903)
         );
  NOR2X1 U17229 ( .A(n27898), .B(n35858), .Y(n27904) );
  AND2XL U17230 ( .A(n23105), .B(n23104), .Y(n28864) );
  NOR2X1 U17231 ( .A(n35858), .B(n33994), .Y(n29062) );
  AOI222XL U17232 ( .A0(n28146), .A1(n28145), .B0(n28146), .B1(conv_2[243]), 
        .C0(n28145), .C1(conv_2[243]), .Y(n28147) );
  NOR2X1 U17233 ( .A(n35858), .B(n28660), .Y(n28664) );
  AND2XL U17234 ( .A(n22901), .B(n22900), .Y(n27971) );
  NOR2X1 U17235 ( .A(n22901), .B(n22900), .Y(n27970) );
  AND2XL U17236 ( .A(n23336), .B(n23335), .Y(n24353) );
  NOR2X1 U17237 ( .A(n23336), .B(n23335), .Y(n24352) );
  NOR2X1 U17238 ( .A(n26509), .B(n35858), .Y(n24015) );
  AOI2BB1XL U17239 ( .A0N(conv_2[18]), .A1N(n27552), .B0(n27551), .Y(n27553)
         );
  NOR2X1 U17240 ( .A(n30195), .B(n35858), .Y(n27554) );
  NAND2XL U17241 ( .A(n34827), .B(n26374), .Y(n21704) );
  AOI22XL U17242 ( .A0(n25289), .A1(conv_3[124]), .B0(n22615), .B1(conv_3[139]), .Y(n19366) );
  AOI22XL U17243 ( .A0(n18658), .A1(conv_3[4]), .B0(n22615), .B1(conv_3[49]), 
        .Y(n18495) );
  AOI2BB2XL U17244 ( .B0(n36245), .B1(n25767), .A0N(n25761), .A1N(n36245), .Y(
        n35108) );
  AOI22XL U17245 ( .A0(n36246), .A1(n20495), .B0(n20490), .B1(n22743), .Y(
        n35104) );
  AND2XL U17246 ( .A(n27626), .B(n27625), .Y(n34092) );
  NOR2X1 U17247 ( .A(n27626), .B(n27625), .Y(n34093) );
  AOI2BB1XL U17248 ( .A0N(conv_3[468]), .A1N(n30184), .B0(n30185), .Y(n19019)
         );
  AND2XL U17249 ( .A(n31695), .B(n31694), .Y(n34072) );
  NOR2X1 U17250 ( .A(n31695), .B(n31694), .Y(n34073) );
  NOR2X1 U17251 ( .A(n31691), .B(n28070), .Y(n26814) );
  NOR2X1 U17252 ( .A(n19108), .B(n31691), .Y(n23223) );
  AOI2BB1XL U17253 ( .A0N(conv_3[228]), .A1N(n29669), .B0(n29670), .Y(n22163)
         );
  NOR2X1 U17254 ( .A(n29136), .B(n31691), .Y(n22164) );
  NOR2X1 U17255 ( .A(n31691), .B(n28660), .Y(n23623) );
  AOI2BB1XL U17256 ( .A0N(conv_3[93]), .A1N(n29637), .B0(n29638), .Y(n22876)
         );
  NOR2X1 U17257 ( .A(n26509), .B(n31691), .Y(n22877) );
  AND2XL U17258 ( .A(n22921), .B(n22920), .Y(n31804) );
  NOR2X1 U17259 ( .A(n22921), .B(n22920), .Y(n31803) );
  AOI222XL U17260 ( .A0(n21702), .A1(n22095), .B0(n21702), .B1(n21701), .C0(
        n22095), .C1(n21700), .Y(n21790) );
  NAND2XL U17261 ( .A(n36246), .B(n25304), .Y(n20185) );
  OAI211XL U17262 ( .A0(n36246), .A1(n22722), .B0(n28528), .C0(n20194), .Y(
        n20195) );
  AOI222XL U17263 ( .A0(n20317), .A1(n20610), .B0(n20317), .B1(n20316), .C0(
        n20610), .C1(n20315), .Y(n20347) );
  NAND2XL U17264 ( .A(n19754), .B(n19753), .Y(n21458) );
  AOI22XL U17265 ( .A0(n36246), .A1(n25298), .B0(n25294), .B1(n22743), .Y(
        n21466) );
  AOI22XL U17266 ( .A0(n36246), .A1(n25304), .B0(n25305), .B1(n22743), .Y(
        n21468) );
  AOI222XL U17267 ( .A0(n20161), .A1(n20039), .B0(n20161), .B1(n20038), .C0(
        n20039), .C1(n20037), .Y(n20097) );
  NOR4BXL U17268 ( .AN(n20036), .B(n20162), .C(n20035), .D(n20034), .Y(n20037)
         );
  AOI222XL U17269 ( .A0(n30647), .A1(n28548), .B0(n30647), .B1(n28547), .C0(
        n28548), .C1(n28546), .Y(n28593) );
  NOR4BBXL U17270 ( .AN(n28545), .BN(n28544), .C(n30646), .D(n28543), .Y(
        n28546) );
  AOI211XL U17271 ( .A0(n34963), .A1(n28412), .B0(n26464), .C0(n26463), .Y(
        n26465) );
  AOI22XL U17272 ( .A0(n28528), .A1(n28560), .B0(n34963), .B1(n28558), .Y(
        n26472) );
  AOI222XL U17273 ( .A0(n26461), .A1(n28617), .B0(n26461), .B1(n26460), .C0(
        n28617), .C1(n26459), .Y(n26490) );
  NOR4XL U17274 ( .A(n28616), .B(n26438), .C(n26437), .D(n26436), .Y(n26460)
         );
  AOI211XL U17275 ( .A0(n34963), .A1(n28583), .B0(n26644), .C0(n26643), .Y(
        n26645) );
  AOI22XL U17276 ( .A0(n34963), .A1(n26632), .B0(n28413), .B1(n16663), .Y(
        n26638) );
  AOI222XL U17277 ( .A0(n26631), .A1(n27979), .B0(n26631), .B1(n26630), .C0(
        n27979), .C1(n26629), .Y(n26663) );
  NOR4XL U17278 ( .A(n27980), .B(n26603), .C(n26602), .D(n26601), .Y(n26630)
         );
  AOI22XL U17279 ( .A0(n25306), .A1(conv_1[75]), .B0(n16662), .B1(conv_1[90]), 
        .Y(n25307) );
  AOI22XL U17280 ( .A0(n36246), .A1(n25305), .B0(n25304), .B1(n21688), .Y(
        n34847) );
  AOI22XL U17281 ( .A0(n25306), .A1(conv_1[315]), .B0(n16673), .B1(conv_1[345]), .Y(n25301) );
  AOI22XL U17282 ( .A0(n25306), .A1(conv_1[375]), .B0(n25299), .B1(conv_1[360]), .Y(n25296) );
  NOR2X1 U17283 ( .A(n29987), .B(n29983), .Y(n29993) );
  AOI2BB1XL U17284 ( .A0N(conv_1[484]), .A1N(n27398), .B0(n27399), .Y(n27220)
         );
  AOI21XL U17285 ( .A0(n27173), .A1(conv_1[473]), .B0(n32887), .Y(n26342) );
  AOI2BB1XL U17286 ( .A0N(conv_1[454]), .A1N(n27392), .B0(n27393), .Y(n27238)
         );
  AOI2BB1XL U17287 ( .A0N(conv_1[439]), .A1N(n27000), .B0(n27001), .Y(n23643)
         );
  AOI2BB1XL U17288 ( .A0N(conv_1[426]), .A1N(intadd_1_n1), .B0(n29328), .Y(
        n29401) );
  NOR2X1 U17289 ( .A(n35501), .B(n35503), .Y(n29402) );
  AOI21XL U17290 ( .A0(n35462), .A1(conv_1[383]), .B0(n35463), .Y(n34336) );
  AOI2BB1XL U17291 ( .A0N(conv_1[364]), .A1N(n30276), .B0(n30277), .Y(n22812)
         );
  NAND2XL U17292 ( .A(n35455), .B(n31365), .Y(n34307) );
  AOI2BB1XL U17293 ( .A0N(conv_1[349]), .A1N(n30282), .B0(n30283), .Y(n24319)
         );
  NOR2X1 U17294 ( .A(n22982), .B(n22981), .Y(n23141) );
  NOR2X1 U17295 ( .A(n33423), .B(n33866), .Y(n19213) );
  NOR2X1 U17296 ( .A(n29197), .B(n29229), .Y(n29280) );
  NOR2X1 U17297 ( .A(n29196), .B(n29195), .Y(n29281) );
  NOR2X1 U17298 ( .A(n33219), .B(n33214), .Y(n24693) );
  NOR2X1 U17299 ( .A(n28601), .B(n28600), .Y(n34300) );
  NAND2X1 U17300 ( .A(n22140), .B(n22139), .Y(n27849) );
  AOI22XL U17301 ( .A0(n26470), .A1(n22850), .B0(n16755), .B1(n22848), .Y(
        n22140) );
  AOI22XL U17302 ( .A0(n28465), .A1(n22818), .B0(n34827), .B1(n22849), .Y(
        n22139) );
  AOI2BB1XL U17303 ( .A0N(conv_1[199]), .A1N(n24168), .B0(n24169), .Y(n23439)
         );
  NAND2XL U17304 ( .A(n35365), .B(n32991), .Y(n34086) );
  AOI2BB1XL U17305 ( .A0N(conv_1[142]), .A1N(n35337), .B0(n32780), .Y(n26765)
         );
  AND2XL U17306 ( .A(n34292), .B(n23650), .Y(n29304) );
  NOR2X1 U17307 ( .A(n31348), .B(n31342), .Y(n34556) );
  OAI21XL U17308 ( .A0(conv_1[109]), .A1(n32880), .B0(n32881), .Y(n24349) );
  AOI2BB1XL U17309 ( .A0N(conv_1[94]), .A1N(n26921), .B0(n26922), .Y(n26514)
         );
  NAND2XL U17310 ( .A(n31337), .B(n26841), .Y(n31335) );
  NOR2X1 U17311 ( .A(conv_1[86]), .B(n26729), .Y(n26737) );
  NOR2X1 U17312 ( .A(n26311), .B(n27088), .Y(n26309) );
  AOI2BB1XL U17313 ( .A0N(conv_1[34]), .A1N(n27036), .B0(n27037), .Y(n25079)
         );
  AOI22XL U17314 ( .A0(n19006), .A1(filter_1[6]), .B0(n19004), .B1(
        filter_1[30]), .Y(n18838) );
  AOI22XL U17315 ( .A0(n19008), .A1(filter_1[42]), .B0(n19007), .B1(
        filter_1[24]), .Y(n18837) );
  OAI2BB1XL U17316 ( .A0N(n19009), .A1N(filter_1[18]), .B0(n18835), .Y(n18839)
         );
  NAND4BX1 U17317 ( .AN(n18729), .B(n18728), .C(n18727), .D(n18726), .Y(n27632) );
  AOI22XL U17318 ( .A0(n19009), .A1(filter_1[23]), .B0(n19006), .B1(
        filter_1[11]), .Y(n18727) );
  AOI22XL U17319 ( .A0(n19004), .A1(filter_1[35]), .B0(filter_1[29]), .B1(
        n19007), .Y(n18728) );
  AOI2BB1XL U17320 ( .A0N(conv_1[19]), .A1N(n27450), .B0(n27451), .Y(n26505)
         );
  INVXL U17321 ( .A(n30672), .Y(n33423) );
  INVXL U17322 ( .A(n21704), .Y(n21756) );
  NAND2XL U17323 ( .A(n34827), .B(n19099), .Y(n21536) );
  OAI22XL U17324 ( .A0(n21033), .A1(n21032), .B0(n21031), .B1(n22052), .Y(
        n21087) );
  NOR4BXL U17325 ( .AN(n21030), .B(n22053), .C(n21029), .D(n21028), .Y(n21031)
         );
  NAND2XL U17326 ( .A(n21831), .B(n25766), .Y(n21960) );
  AOI22XL U17327 ( .A0(n25306), .A1(conv_2[345]), .B0(n18810), .B1(conv_2[360]), .Y(n20741) );
  AOI22XL U17328 ( .A0(n25299), .A1(conv_2[330]), .B0(n22615), .B1(conv_2[375]), .Y(n20740) );
  AOI222XL U17329 ( .A0(n21975), .A1(n22189), .B0(n21975), .B1(n21974), .C0(
        n22189), .C1(n21973), .Y(n22046) );
  NOR4XL U17330 ( .A(n22188), .B(n21972), .C(n21971), .D(n21938), .Y(n21974)
         );
  AOI211XL U17331 ( .A0(n34963), .A1(n25651), .B0(n25045), .C0(n25044), .Y(
        n25047) );
  NAND2XL U17332 ( .A(n34963), .B(n25643), .Y(n25040) );
  NOR2X1 U17333 ( .A(n25636), .B(n16721), .Y(n25039) );
  AOI222XL U17334 ( .A0(n25029), .A1(n25443), .B0(n25029), .B1(n25028), .C0(
        n25443), .C1(n25027), .Y(n25058) );
  NOR4XL U17335 ( .A(n25444), .B(n25024), .C(n25023), .D(n25022), .Y(n25028)
         );
  AOI222XL U17336 ( .A0(n26349), .A1(n25198), .B0(n26349), .B1(n25197), .C0(
        n25198), .C1(n25196), .Y(n25227) );
  NOR2X1 U17337 ( .A(n35261), .B(n28391), .Y(n28595) );
  AOI22XL U17338 ( .A0(n34963), .A1(n34930), .B0(n16670), .B1(n25100), .Y(
        n24048) );
  OAI2BB2XL U17339 ( .B0(n24111), .B1(n24110), .A0N(pool[59]), .A1N(n24109), 
        .Y(n24132) );
  AOI22XL U17340 ( .A0(n34963), .A1(n25632), .B0(n16670), .B1(n25635), .Y(
        n24787) );
  AOI211XL U17341 ( .A0(n34963), .A1(n25628), .B0(n24780), .C0(n24779), .Y(
        n24781) );
  AOI222XL U17342 ( .A0(n24777), .A1(n26151), .B0(n24777), .B1(n24776), .C0(
        n26151), .C1(n24775), .Y(n24804) );
  NOR4XL U17343 ( .A(n26150), .B(n24756), .C(n24755), .D(n24754), .Y(n24776)
         );
  AOI22XL U17344 ( .A0(n36246), .A1(n24043), .B0(n24042), .B1(n21688), .Y(
        n34931) );
  OAI222XL U17345 ( .A0(n24041), .A1(n22612), .B0(n36246), .B1(n24040), .C0(
        n34456), .C1(n24039), .Y(n34932) );
  AOI222XL U17346 ( .A0(n25617), .A1(n27372), .B0(n25617), .B1(n25616), .C0(
        n27372), .C1(n25615), .Y(n25671) );
  NOR4XL U17347 ( .A(n27371), .B(n25555), .C(n25554), .D(n25612), .Y(n25616)
         );
  AOI2BB1XL U17348 ( .A0N(conv_2[517]), .A1N(n27787), .B0(n28706), .Y(n27781)
         );
  NOR2X1 U17349 ( .A(n27792), .B(n27788), .Y(n27782) );
  AOI2BB1XL U17350 ( .A0N(conv_2[514]), .A1N(n28971), .B0(n28972), .Y(n27771)
         );
  NOR2X1 U17351 ( .A(n30911), .B(n30910), .Y(n36074) );
  AOI2BB1XL U17352 ( .A0N(conv_2[484]), .A1N(n28983), .B0(n28984), .Y(n27741)
         );
  OR2XL U17353 ( .A(n27943), .B(n27881), .Y(n34171) );
  NOR2X1 U17354 ( .A(n27881), .B(n30900), .Y(n34172) );
  OR2XL U17355 ( .A(n27943), .B(n27867), .Y(n33892) );
  INVXL U17356 ( .A(n34173), .Y(n27943) );
  OAI21XL U17357 ( .A0(conv_2[455]), .A1(n30876), .B0(n33611), .Y(n30877) );
  INVXL U17358 ( .A(n29046), .Y(n35858) );
  AOI2BB1XL U17359 ( .A0N(conv_2[440]), .A1N(n28943), .B0(n28937), .Y(n36059)
         );
  NOR2X1 U17360 ( .A(n28942), .B(n28947), .Y(n36060) );
  AOI2BB1XL U17361 ( .A0N(conv_2[439]), .A1N(n29028), .B0(n29029), .Y(n27905)
         );
  INVXL U17362 ( .A(n34224), .Y(n27898) );
  NAND2XL U17363 ( .A(n36067), .B(n27923), .Y(n30962) );
  AOI2BB1XL U17364 ( .A0N(conv_2[424]), .A1N(n29016), .B0(n29017), .Y(n28133)
         );
  AOI2BB1XL U17365 ( .A0N(conv_2[379]), .A1N(n29010), .B0(n29011), .Y(n23079)
         );
  NAND2XL U17366 ( .A(n18741), .B(n18740), .Y(n22802) );
  NOR2X1 U17367 ( .A(n29518), .B(n29522), .Y(n29525) );
  OR2XL U17368 ( .A(n33925), .B(n33924), .Y(n33926) );
  NOR2X1 U17369 ( .A(n33989), .B(n34418), .Y(n23096) );
  AND2XL U17370 ( .A(n35982), .B(n23106), .Y(n28050) );
  AOI2BB1XL U17371 ( .A0N(conv_2[304]), .A1N(n28870), .B0(n28871), .Y(n19114)
         );
  AOI2BB1XL U17372 ( .A0N(conv_2[289]), .A1N(n29034), .B0(n29035), .Y(n28091)
         );
  NAND2XL U17373 ( .A(n18803), .B(n18802), .Y(n22817) );
  AOI222XL U17374 ( .A0(n29408), .A1(n29409), .B0(n29408), .B1(conv_2[259]), 
        .C0(n29409), .C1(conv_2[259]), .Y(n19043) );
  AND2XL U17375 ( .A(n33770), .B(n28665), .Y(n29915) );
  AOI2BB1XL U17376 ( .A0N(conv_2[184]), .A1N(n29022), .B0(n29023), .Y(n28655)
         );
  AOI2BB1XL U17377 ( .A0N(conv_2[172]), .A1N(n29846), .B0(n33974), .Y(n29852)
         );
  AOI2BB1XL U17378 ( .A0N(conv_2[169]), .A1N(n29833), .B0(n29832), .Y(n29834)
         );
  NOR2X1 U17379 ( .A(n34627), .B(n28631), .Y(n34624) );
  NOR2X1 U17380 ( .A(n23115), .B(n23114), .Y(n23369) );
  AND2XL U17381 ( .A(n23115), .B(n23114), .Y(n23370) );
  NAND2XL U17382 ( .A(n18962), .B(n18961), .Y(n22936) );
  AOI22XL U17383 ( .A0(n22370), .A1(n23240), .B0(n21100), .B1(n19051), .Y(
        n18962) );
  AOI22XL U17384 ( .A0(n22362), .A1(n19052), .B0(n22369), .B1(n23239), .Y(
        n18961) );
  NAND2XL U17385 ( .A(n34626), .B(n24531), .Y(n33947) );
  OAI2BB1XL U17386 ( .A0N(conv_2[160]), .A1N(n34624), .B0(n34623), .Y(n33946)
         );
  AOI2BB1XL U17387 ( .A0N(conv_2[139]), .A1N(n27971), .B0(n27970), .Y(n27972)
         );
  AOI2BB1XL U17388 ( .A0N(conv_2[124]), .A1N(n24353), .B0(n24352), .Y(n24354)
         );
  OAI2BB1XL U17389 ( .A0N(conv_2[115]), .A1N(n30149), .B0(n35884), .Y(n34642)
         );
  NAND2XL U17390 ( .A(n30225), .B(n30204), .Y(n30938) );
  INVXL U17391 ( .A(n30940), .Y(n30225) );
  AOI2BB1XL U17392 ( .A0N(conv_2[79]), .A1N(n28741), .B0(n28740), .Y(n28742)
         );
  AOI21XL U17393 ( .A0(conv_2[70]), .A1(n30126), .B0(n33735), .Y(n30241) );
  NOR2X1 U17394 ( .A(n30120), .B(n30119), .Y(n30973) );
  NOR2X1 U17395 ( .A(n33586), .B(n35862), .Y(n29618) );
  AOI22XL U17396 ( .A0(n19009), .A1(filter_2[23]), .B0(n19008), .B1(
        filter_2[47]), .Y(n18899) );
  AOI22XL U17397 ( .A0(n19006), .A1(filter_2[11]), .B0(n19007), .B1(
        filter_2[29]), .Y(n18900) );
  AOI2BB2XL U17398 ( .B0(n16665), .B1(n34955), .A0N(n34959), .A1N(n28575), .Y(
        n21115) );
  AOI222XL U17399 ( .A0(n21380), .A1(n22108), .B0(n21380), .B1(n21379), .C0(
        n22108), .C1(n21378), .Y(n21454) );
  AOI22XL U17400 ( .A0(n25289), .A1(conv_3[360]), .B0(n18240), .B1(conv_3[375]), .Y(n19256) );
  AOI22XL U17401 ( .A0(n25289), .A1(conv_3[120]), .B0(n22615), .B1(conv_3[135]), .Y(n19255) );
  AOI22XL U17402 ( .A0(n25289), .A1(conv_3[60]), .B0(n22690), .B1(conv_3[30]), 
        .Y(n19261) );
  AOI22XL U17403 ( .A0(n25289), .A1(conv_3[300]), .B0(n22615), .B1(conv_3[315]), .Y(n19264) );
  INVXL U17404 ( .A(n21830), .Y(n21831) );
  AOI22XL U17405 ( .A0(n36246), .A1(n22226), .B0(n22227), .B1(n22713), .Y(
        n34953) );
  INVXL U17406 ( .A(n21960), .Y(n34950) );
  AOI22XL U17407 ( .A0(n36244), .A1(n35169), .B0(n34963), .B1(n28265), .Y(
        n26168) );
  AOI211XL U17408 ( .A0(n34963), .A1(n35180), .B0(n26282), .C0(n26281), .Y(
        n26284) );
  NOR2X1 U17409 ( .A(n35182), .B(n26274), .Y(n26282) );
  AOI222XL U17410 ( .A0(n26258), .A1(n27066), .B0(n26258), .B1(n26257), .C0(
        n27066), .C1(n26256), .Y(n26292) );
  NOR4XL U17411 ( .A(n26252), .B(n26253), .C(n27067), .D(n26236), .Y(n26257)
         );
  INVXL U17412 ( .A(n25337), .Y(n25402) );
  AOI22XL U17413 ( .A0(n34963), .A1(n28365), .B0(n16670), .B1(n35185), .Y(
        n18687) );
  AOI22XL U17414 ( .A0(n34963), .A1(n28373), .B0(n28324), .B1(n35193), .Y(
        n18704) );
  NAND2XL U17415 ( .A(n19767), .B(n26274), .Y(n26451) );
  NOR2X1 U17416 ( .A(n22847), .B(n25766), .Y(n28304) );
  NOR4XL U17417 ( .A(n28385), .B(n28384), .C(n28383), .D(n28382), .Y(n28386)
         );
  NAND2XL U17418 ( .A(n22234), .B(n22233), .Y(n28293) );
  AOI22XL U17419 ( .A0(n25306), .A1(conv_3[315]), .B0(n22615), .B1(conv_3[345]), .Y(n22233) );
  NAND2XL U17420 ( .A(n22241), .B(n22240), .Y(n34986) );
  NAND2X1 U17421 ( .A(n23053), .B(n26285), .Y(n35231) );
  NAND2XL U17422 ( .A(n22229), .B(n22228), .Y(n35232) );
  AOI22XL U17423 ( .A0(n18658), .A1(conv_3[360]), .B0(n22615), .B1(conv_3[405]), .Y(n22236) );
  AOI22XL U17424 ( .A0(n36246), .A1(n22227), .B0(n22226), .B1(n21688), .Y(
        n35230) );
  AOI222XL U17425 ( .A0(n26708), .A1(n25785), .B0(n26708), .B1(n25784), .C0(
        n25785), .C1(n25783), .Y(n25807) );
  NOR4BBXL U17426 ( .AN(n25782), .BN(n25781), .C(n25780), .D(n26707), .Y(
        n25783) );
  AOI2BB1XL U17427 ( .A0N(conv_3[499]), .A1N(n34092), .B0(n34093), .Y(n27627)
         );
  AOI2BB1XL U17428 ( .A0N(conv_3[469]), .A1N(n22190), .B0(n22191), .Y(n19021)
         );
  AOI222XL U17429 ( .A0(n24260), .A1(n24261), .B0(n24260), .B1(conv_3[454]), 
        .C0(n24261), .C1(conv_3[454]), .Y(n19062) );
  AOI22XL U17430 ( .A0(n22369), .A1(n19051), .B0(n22370), .B1(n19050), .Y(
        n22800) );
  AOI2BB1XL U17431 ( .A0N(conv_3[439]), .A1N(n31926), .B0(n31925), .Y(n31927)
         );
  NAND2XL U17432 ( .A(n22206), .B(n22205), .Y(n23090) );
  NOR2X1 U17433 ( .A(conv_3[431]), .B(n32157), .Y(n32581) );
  AOI2BB1XL U17434 ( .A0N(conv_3[429]), .A1N(n35773), .B0(n35775), .Y(n31726)
         );
  AOI2BB1XL U17435 ( .A0N(conv_3[424]), .A1N(n34072), .B0(n34073), .Y(n31696)
         );
  NAND2XL U17436 ( .A(n18761), .B(n18760), .Y(n22937) );
  AOI22XL U17437 ( .A0(n22370), .A1(n23242), .B0(n21100), .B1(n23244), .Y(
        n18760) );
  AOI22XL U17438 ( .A0(n22362), .A1(n23241), .B0(n22369), .B1(n23243), .Y(
        n18761) );
  INVXL U17439 ( .A(n32557), .Y(n32558) );
  AOI2BB1XL U17440 ( .A0N(conv_3[394]), .A1N(n32019), .B0(n32018), .Y(n32020)
         );
  OR2X1 U17441 ( .A(n32200), .B(n32199), .Y(n34162) );
  NOR2X1 U17442 ( .A(n32199), .B(n32198), .Y(n34163) );
  AOI2BB1XL U17443 ( .A0N(conv_3[364]), .A1N(n31626), .B0(n31625), .Y(n31627)
         );
  NOR2X1 U17444 ( .A(conv_3[356]), .B(n32128), .Y(n32131) );
  AOI2BB1XL U17445 ( .A0N(conv_3[304]), .A1N(n31405), .B0(n31404), .Y(n31406)
         );
  AND2XL U17446 ( .A(n23066), .B(n23065), .Y(n23666) );
  NOR2X1 U17447 ( .A(n23066), .B(n23065), .Y(n23667) );
  AOI2BB1XL U17448 ( .A0N(conv_3[276]), .A1N(n31744), .B0(n32599), .Y(n31750)
         );
  AOI2BB1XL U17449 ( .A0N(conv_3[244]), .A1N(n28797), .B0(n28796), .Y(n28798)
         );
  OAI21XL U17450 ( .A0(conv_3[235]), .A1(n31060), .B0(n35673), .Y(n33314) );
  AOI2BB1XL U17451 ( .A0N(conv_3[229]), .A1N(n26153), .B0(n26152), .Y(n26154)
         );
  AOI2BB1XL U17452 ( .A0N(conv_3[214]), .A1N(n26525), .B0(n26524), .Y(n26526)
         );
  OAI21XL U17453 ( .A0(conv_3[199]), .A1(n24474), .B0(n24473), .Y(n24475) );
  INVX2 U17454 ( .A(n27849), .Y(n27848) );
  AOI2BB1XL U17455 ( .A0N(conv_3[184]), .A1N(n26316), .B0(n26315), .Y(n26317)
         );
  NOR2X1 U17456 ( .A(n31561), .B(n31560), .Y(n31562) );
  INVXL U17457 ( .A(n35639), .Y(n32221) );
  AOI2BB1XL U17458 ( .A0N(conv_3[154]), .A1N(n29746), .B0(n29745), .Y(n29747)
         );
  OR2XL U17459 ( .A(n32789), .B(n23778), .Y(n34395) );
  AOI2BB1XL U17460 ( .A0N(conv_3[124]), .A1N(n28950), .B0(n28949), .Y(n28951)
         );
  AOI2BB1XL U17461 ( .A0N(conv_3[94]), .A1N(n31667), .B0(n31666), .Y(n31668)
         );
  NAND2XL U17462 ( .A(n34186), .B(n32116), .Y(n34188) );
  AOI22XL U17463 ( .A0(n19008), .A1(filter_3[47]), .B0(n19004), .B1(
        filter_3[35]), .Y(n18979) );
  AOI22XL U17464 ( .A0(n19006), .A1(filter_3[11]), .B0(n19007), .B1(
        filter_3[29]), .Y(n18978) );
  AOI2BB1XL U17465 ( .A0N(conv_3[79]), .A1N(n31804), .B0(n31803), .Y(n31805)
         );
  NAND4BX2 U17466 ( .AN(n19002), .B(n19001), .C(n19000), .D(n18999), .Y(n29678) );
  AOI22XL U17467 ( .A0(n19009), .A1(filter_3[18]), .B0(n19004), .B1(
        filter_3[30]), .Y(n19000) );
  AOI22XL U17468 ( .A0(n19007), .A1(filter_3[24]), .B0(n19005), .B1(
        filter_3[12]), .Y(n18999) );
  INVXL U17469 ( .A(n24467), .Y(n31691) );
  NOR2X1 U17470 ( .A(n20178), .B(n20172), .Y(n20170) );
  NAND2XL U17471 ( .A(n20165), .B(n26846), .Y(n30350) );
  NAND2X1 U17472 ( .A(counter[1]), .B(counter[0]), .Y(n19245) );
  NAND2XL U17473 ( .A(n18175), .B(n18176), .Y(n18189) );
  NOR3X1 U17474 ( .A(n18158), .B(n19245), .C(n18157), .Y(n18185) );
  AOI21XL U17475 ( .A0(n20165), .A1(n18159), .B0(cs[2]), .Y(n18177) );
  NAND2XL U17476 ( .A(counter[2]), .B(n17988), .Y(n18174) );
  NAND2XL U17477 ( .A(n18191), .B(cs[0]), .Y(n18173) );
  NAND2XL U17478 ( .A(n29676), .B(weight_1_bias_1[5]), .Y(n33077) );
  NAND2XL U17479 ( .A(n29676), .B(weight_1_bias_2[5]), .Y(n33564) );
  NAND2XL U17480 ( .A(n29676), .B(weight_1_bias_3[5]), .Y(n33412) );
  NAND2XL U17481 ( .A(weight_2_bias_2[5]), .B(n20614), .Y(n33350) );
  NOR2X1 U17482 ( .A(n35272), .B(n34770), .Y(n33401) );
  NOR2X1 U17483 ( .A(n24554), .B(n24552), .Y(n24550) );
  NOR2X1 U17484 ( .A(n30536), .B(n28762), .Y(n27478) );
  NOR2X1 U17485 ( .A(n23744), .B(n23746), .Y(n23742) );
  AND2XL U17486 ( .A(n24909), .B(n22217), .Y(n30460) );
  NOR2X1 U17487 ( .A(n30486), .B(n30485), .Y(n30488) );
  ADDFXL U17488 ( .A(conv_1[362]), .B(n24232), .CI(n24231), .CO(n28965), .S(
        n24234) );
  NOR2X1 U17489 ( .A(n33403), .B(n23504), .Y(n24232) );
  OAI2BB2XL U17490 ( .B0(n35272), .B1(n30057), .A0N(n30132), .A1N(conv_1[361]), 
        .Y(n24231) );
  OAI2BB1XL U17491 ( .A0N(n33134), .A1N(n29676), .B0(n25246), .Y(n24233) );
  ADDFHX1 U17492 ( .A(conv_2[512]), .B(n27766), .CI(n27765), .CO(n29645), .S(
        n23566) );
  OAI31XL U17493 ( .A0(n35853), .A1(n27644), .A2(n23719), .B0(n23718), .Y(
        n30015) );
  OAI2BB1XL U17494 ( .A0N(n30254), .A1N(n29676), .B0(n24279), .Y(n23575) );
  ADDFXL U17495 ( .A(conv_3[377]), .B(n24247), .CI(n24246), .CO(n19191), .S(
        n24248) );
  NOR2X1 U17496 ( .A(n18997), .B(n27532), .Y(n24247) );
  ADDFXL U17497 ( .A(conv_3[362]), .B(n23562), .CI(n23561), .CO(n23505), .S(
        n23563) );
  AOI2BB1XL U17498 ( .A0N(conv_3[361]), .A1N(n30562), .B0(n30563), .Y(n23561)
         );
  ADDFXL U17499 ( .A(conv_3[272]), .B(n33024), .CI(n33023), .CO(n23493), .S(
        n33025) );
  NOR2XL U17500 ( .A(n18997), .B(n33994), .Y(n33024) );
  NOR2X1 U17501 ( .A(n23423), .B(n23422), .Y(n29542) );
  ADDFXL U17502 ( .A(conv_1[393]), .B(n27634), .CI(n27633), .CO(n27635), .S(
        n23021) );
  NOR2X1 U17503 ( .A(n35498), .B(n32016), .Y(n27634) );
  OAI2BB1XL U17504 ( .A0N(conv_1[317]), .A1N(n30494), .B0(n22274), .Y(n22437)
         );
  OAI2BB1XL U17505 ( .A0N(n23162), .A1N(n29676), .B0(n24673), .Y(n24288) );
  AND2XL U17506 ( .A(n23468), .B(n23467), .Y(n24690) );
  ADDFXL U17507 ( .A(conv_1[213]), .B(n24292), .CI(n24291), .CO(n23999), .S(
        n24294) );
  NOR2X1 U17508 ( .A(n35498), .B(n28660), .Y(n24292) );
  OAI2BB1XL U17509 ( .A0N(n28606), .A1N(n29676), .B0(n24673), .Y(n24293) );
  NOR2X1 U17510 ( .A(n35498), .B(n23296), .Y(n24283) );
  OAI2BB1XL U17511 ( .A0N(n31341), .A1N(n29676), .B0(n24673), .Y(n26515) );
  NOR2XL U17512 ( .A(n35498), .B(n31418), .Y(n26140) );
  AOI2BB1XL U17513 ( .A0N(conv_1[62]), .A1N(n26990), .B0(n26991), .Y(n26139)
         );
  NOR2X1 U17514 ( .A(n27902), .B(n27901), .Y(n29553) );
  AND2XL U17515 ( .A(n24449), .B(n24448), .Y(n29565) );
  NOR2X1 U17516 ( .A(n24449), .B(n24448), .Y(n29566) );
  ADDFXL U17517 ( .A(conv_2[348]), .B(n23713), .CI(n23712), .CO(n24193), .S(
        n23714) );
  ADDFXL U17518 ( .A(conv_2[333]), .B(n24302), .CI(n24301), .CO(n23868), .S(
        n24304) );
  NOR2X1 U17519 ( .A(n35856), .B(n33994), .Y(n23703) );
  ADDFXL U17520 ( .A(conv_2[213]), .B(n28662), .CI(n28661), .CO(n28663), .S(
        n23710) );
  ADDFXL U17521 ( .A(conv_2[93]), .B(n23032), .CI(n23031), .CO(n24016), .S(
        n23034) );
  OAI2BB1XL U17522 ( .A0N(n30232), .A1N(n29676), .B0(n24279), .Y(n23033) );
  NOR2X1 U17523 ( .A(n23795), .B(n23794), .Y(n27701) );
  NOR2X1 U17524 ( .A(n23581), .B(n23580), .Y(n27552) );
  AND2XL U17525 ( .A(n23581), .B(n23580), .Y(n27551) );
  ADDFXL U17526 ( .A(conv_3[513]), .B(n23739), .CI(n23738), .CO(n23260), .S(
        n23740) );
  NOR2XL U17527 ( .A(n29426), .B(n27764), .Y(n23739) );
  ADDFXL U17528 ( .A(conv_3[483]), .B(n23515), .CI(n23514), .CO(n23516), .S(
        n23062) );
  NOR2X1 U17529 ( .A(n27735), .B(n29426), .Y(n23515) );
  NOR2X1 U17530 ( .A(n19018), .B(n19017), .Y(n30184) );
  AND2XL U17531 ( .A(n19018), .B(n19017), .Y(n30185) );
  NOR2X1 U17532 ( .A(n29684), .B(n29683), .Y(n31693) );
  AND2XL U17533 ( .A(n29684), .B(n29683), .Y(n31692) );
  NOR2X1 U17534 ( .A(n29426), .B(n28070), .Y(n24327) );
  AOI2BB1XL U17535 ( .A0N(conv_3[407]), .A1N(n30543), .B0(n30544), .Y(n24326)
         );
  ADDFXL U17536 ( .A(conv_3[348]), .B(n26716), .CI(n26715), .CO(n31391), .S(
        n24335) );
  AND2XL U17537 ( .A(n22113), .B(n22112), .Y(n29414) );
  NOR2X1 U17538 ( .A(n22113), .B(n22112), .Y(n29415) );
  NOR2X1 U17539 ( .A(n22162), .B(n22161), .Y(n29669) );
  AND2XL U17540 ( .A(n22162), .B(n22161), .Y(n29670) );
  ADDFXL U17541 ( .A(conv_3[213]), .B(n24323), .CI(n24322), .CO(n23622), .S(
        n24324) );
  NOR2X1 U17542 ( .A(n29426), .B(n28660), .Y(n24323) );
  NOR2X1 U17543 ( .A(n22875), .B(n22874), .Y(n29637) );
  AND2XL U17544 ( .A(n22875), .B(n22874), .Y(n29638) );
  OAI2BB1XL U17545 ( .A0N(n32156), .A1N(n29676), .B0(n25246), .Y(n23731) );
  NOR2X1 U17546 ( .A(n30195), .B(n29426), .Y(n29978) );
  NOR2X1 U17547 ( .A(n29426), .B(n35857), .Y(n24331) );
  INVXL U17548 ( .A(n34815), .Y(n34813) );
  INVXL U17549 ( .A(n34844), .Y(n34840) );
  INVXL U17550 ( .A(n34800), .Y(n34798) );
  INVXL U17551 ( .A(n34821), .Y(n34817) );
  INVXL U17552 ( .A(n34806), .Y(n34802) );
  INVXL U17553 ( .A(n34810), .Y(n34808) );
  AND2XL U17554 ( .A(n27219), .B(n27218), .Y(n27398) );
  AND2XL U17555 ( .A(n18854), .B(n18853), .Y(n27006) );
  NOR2X1 U17556 ( .A(n18854), .B(n18853), .Y(n27007) );
  AND2XL U17557 ( .A(n27636), .B(n27635), .Y(n30759) );
  NOR2X1 U17558 ( .A(n27636), .B(n27635), .Y(n30760) );
  OAI2BB1XL U17559 ( .A0N(n28828), .A1N(n29676), .B0(n24279), .Y(n24242) );
  NOR2X1 U17560 ( .A(n35500), .B(n19108), .Y(n22946) );
  AOI2BB1XL U17561 ( .A0N(conv_1[303]), .A1N(n24224), .B0(n24225), .Y(n22945)
         );
  AND2XL U17562 ( .A(n22298), .B(n22297), .Y(n23909) );
  NOR2X1 U17563 ( .A(n35500), .B(n33020), .Y(n22953) );
  AND2XL U17564 ( .A(n26504), .B(n26503), .Y(n27450) );
  NOR2X1 U17565 ( .A(n35500), .B(n35857), .Y(intadd_2_B_2_) );
  INVXL U17566 ( .A(n34890), .Y(n34888) );
  INVXL U17567 ( .A(n34871), .Y(n34872) );
  INVXL U17568 ( .A(n34866), .Y(n34864) );
  INVXL U17569 ( .A(n34896), .Y(n34892) );
  INVXL U17570 ( .A(n34884), .Y(n34885) );
  INVXL U17571 ( .A(n34901), .Y(n34897) );
  AND2XL U17572 ( .A(n27904), .B(n27903), .Y(n29028) );
  NOR2X1 U17573 ( .A(n27904), .B(n27903), .Y(n29029) );
  AND2XL U17574 ( .A(n28132), .B(n28131), .Y(n29016) );
  NOR2X1 U17575 ( .A(n28132), .B(n28131), .Y(n29017) );
  AND2XL U17576 ( .A(n28664), .B(n28663), .Y(n28876) );
  AND2XL U17577 ( .A(n27554), .B(n27553), .Y(n29713) );
  NOR2X1 U17578 ( .A(n35858), .B(n35857), .Y(intadd_0_B_2_) );
  INVXL U17579 ( .A(n35014), .Y(n35015) );
  INVXL U17580 ( .A(n35026), .Y(n35027) );
  INVXL U17581 ( .A(n34945), .Y(n34948) );
  INVXL U17582 ( .A(n24569), .Y(n35018) );
  NOR2X1 U17583 ( .A(n34093), .B(n34092), .Y(n34095) );
  AND2XL U17584 ( .A(n19020), .B(n19019), .Y(n22190) );
  NOR2X1 U17585 ( .A(n19020), .B(n19019), .Y(n22191) );
  NOR2X1 U17586 ( .A(n34073), .B(n34072), .Y(n34075) );
  AND2XL U17587 ( .A(n23223), .B(n23222), .Y(n31405) );
  AND2XL U17588 ( .A(n24026), .B(n24025), .Y(n28797) );
  NOR2X1 U17589 ( .A(n24026), .B(n24025), .Y(n28796) );
  AND2XL U17590 ( .A(n22164), .B(n22163), .Y(n26153) );
  AND2XL U17591 ( .A(n23623), .B(n23622), .Y(n26525) );
  NOR2X1 U17592 ( .A(n23623), .B(n23622), .Y(n26524) );
  AND2XL U17593 ( .A(n22877), .B(n22876), .Y(n31667) );
  AOI2BB1XL U17594 ( .A0N(conv_1[532]), .A1N(n29209), .B0(n29236), .Y(n29234)
         );
  INVXL U17595 ( .A(n29216), .Y(n29236) );
  MXI2XL U17596 ( .A(n29216), .B(n29236), .S0(n23696), .Y(n23698) );
  AOI22XL U17597 ( .A0(n25289), .A1(conv_1[30]), .B0(n18240), .B1(conv_1[45]), 
        .Y(n25291) );
  OAI2BB1XL U17598 ( .A0N(n25434), .A1N(n28391), .B0(n35227), .Y(n34795) );
  AOI222XL U17599 ( .A0(n25433), .A1(n25432), .B0(n25433), .B1(n25431), .C0(
        n25432), .C1(n25430), .Y(n25434) );
  AOI211XL U17600 ( .A0(n26263), .A1(n26632), .B0(n25317), .C0(n25316), .Y(
        n25433) );
  OAI21XL U17601 ( .A0(n35229), .A1(n24665), .B0(n35227), .Y(n34860) );
  AOI222XL U17602 ( .A0(n24664), .A1(n24663), .B0(n24664), .B1(n24662), .C0(
        n24663), .C1(n24661), .Y(n24665) );
  OAI211XL U17603 ( .A0(n35135), .A1(n26639), .B0(n24638), .C0(n24637), .Y(
        n24663) );
  OAI21XL U17604 ( .A0(n35229), .A1(n22795), .B0(n35227), .Y(n34839) );
  AOI222XL U17605 ( .A0(n22794), .A1(n22793), .B0(n22794), .B1(n22792), .C0(
        n22793), .C1(n22791), .Y(n22795) );
  AOI21XL U17606 ( .A0(n28005), .A1(n29676), .B0(n18856), .Y(n33432) );
  AOI21XL U17607 ( .A0(n29250), .A1(n29676), .B0(n18856), .Y(n35547) );
  NOR2X1 U17608 ( .A(n27131), .B(n27119), .Y(n23428) );
  AOI2BB1XL U17609 ( .A0N(conv_1[499]), .A1N(n30695), .B0(n30696), .Y(n23662)
         );
  OAI2BB1XL U17610 ( .A0N(n27190), .A1N(n29676), .B0(n25246), .Y(n23663) );
  AOI22XL U17611 ( .A0(n23055), .A1(n22151), .B0(n34906), .B1(n22266), .Y(
        n18896) );
  AOI22XL U17612 ( .A0(n25766), .A1(n22447), .B0(n34921), .B1(n22152), .Y(
        n18895) );
  INVXL U17613 ( .A(n35534), .Y(n35541) );
  AND2XL U17614 ( .A(n35541), .B(n27220), .Y(n29971) );
  AOI21XL U17615 ( .A0(n33358), .A1(n29676), .B0(n18856), .Y(n35544) );
  AOI21XL U17616 ( .A0(n28738), .A1(n29676), .B0(n18856), .Y(n33506) );
  AOI2BB1XL U17617 ( .A0N(conv_1[458]), .A1N(n30036), .B0(n30051), .Y(n30031)
         );
  AOI21XL U17618 ( .A0(conv_1[458]), .A1(n30037), .B0(n30044), .Y(n30030) );
  AOI2BB1XL U17619 ( .A0N(conv_1[457]), .A1N(n30049), .B0(n30051), .Y(n30036)
         );
  NOR2X1 U17620 ( .A(n30055), .B(n30050), .Y(n30037) );
  AND2XL U17621 ( .A(n30044), .B(n27238), .Y(n27244) );
  AOI21XL U17622 ( .A0(n28754), .A1(n29676), .B0(n18856), .Y(n30056) );
  OAI2BB1XL U17623 ( .A0N(n27197), .A1N(n29676), .B0(n25246), .Y(n35517) );
  AND2XL U17624 ( .A(n35515), .B(n23643), .Y(n27166) );
  INVXL U17625 ( .A(n35517), .Y(n35520) );
  AOI2BB1XL U17626 ( .A0N(conv_1[427]), .A1N(n29401), .B0(n29328), .Y(n27583)
         );
  INVXL U17627 ( .A(intadd_1_B_2_), .Y(n29328) );
  NOR2X1 U17628 ( .A(conv_1[428]), .B(n27583), .Y(n27582) );
  OAI2BB1XL U17629 ( .A0N(n29334), .A1N(n29676), .B0(n25246), .Y(n35510) );
  AOI2BB1XL U17630 ( .A0N(conv_1[415]), .A1N(n29298), .B0(n29299), .Y(n32687)
         );
  NOR2X1 U17631 ( .A(n27596), .B(n27597), .Y(n33387) );
  OAI2BB1XL U17632 ( .A0N(n34675), .A1N(n29676), .B0(n25246), .Y(n35495) );
  INVXL U17633 ( .A(n35495), .Y(n35487) );
  INVXL U17634 ( .A(n35493), .Y(n34775) );
  NOR2X1 U17635 ( .A(n33652), .B(n35471), .Y(n35476) );
  NOR2X1 U17636 ( .A(conv_1[400]), .B(n33651), .Y(n33652) );
  NOR2X1 U17637 ( .A(n35473), .B(n35470), .Y(n33653) );
  AOI2BB1XL U17638 ( .A0N(conv_1[399]), .A1N(n35469), .B0(n35471), .Y(n33651)
         );
  OAI2BB1XL U17639 ( .A0N(n33273), .A1N(n29676), .B0(n25246), .Y(n33649) );
  AOI2BB1XL U17640 ( .A0N(conv_1[398]), .A1N(n31280), .B0(n35471), .Y(n35469)
         );
  NAND2XL U17641 ( .A(n27632), .B(n27990), .Y(n35471) );
  INVXL U17642 ( .A(n35471), .Y(n33654) );
  AND2XL U17643 ( .A(n33654), .B(n27637), .Y(n29275) );
  NOR2X1 U17644 ( .A(n33654), .B(n27637), .Y(n29274) );
  OAI2BB1XL U17645 ( .A0N(n33152), .A1N(n29676), .B0(n25246), .Y(n22976) );
  INVXL U17646 ( .A(n22976), .Y(n35466) );
  AOI2BB1XL U17647 ( .A0N(conv_1[369]), .A1N(n23151), .B0(n31363), .Y(n31364)
         );
  NOR2X1 U17648 ( .A(n23150), .B(n23149), .Y(n31362) );
  AOI2BB1XL U17649 ( .A0N(conv_1[368]), .A1N(n35453), .B0(n31363), .Y(n23151)
         );
  NAND2XL U17650 ( .A(n27632), .B(n34502), .Y(n31363) );
  INVXL U17651 ( .A(n31363), .Y(n35455) );
  AND2XL U17652 ( .A(n35455), .B(n22812), .Y(n22838) );
  INVXL U17653 ( .A(n24233), .Y(n35458) );
  AND2XL U17654 ( .A(n35441), .B(n24319), .Y(n26363) );
  INVXL U17655 ( .A(n34763), .Y(n35447) );
  OAI2BB1XL U17656 ( .A0N(n28820), .A1N(n29676), .B0(n24279), .Y(n34763) );
  INVXL U17657 ( .A(n24242), .Y(n35437) );
  AOI2BB1XL U17658 ( .A0N(conv_1[324]), .A1N(n23309), .B0(n23310), .Y(n22926)
         );
  AOI2BB1XL U17659 ( .A0N(conv_1[323]), .A1N(n23315), .B0(n29382), .Y(n23309)
         );
  OAI2BB1XL U17660 ( .A0N(n22930), .A1N(n29676), .B0(n24279), .Y(n25268) );
  INVXL U17661 ( .A(n25268), .Y(n34263) );
  OAI2BB1XL U17662 ( .A0N(n24814), .A1N(n29676), .B0(n24279), .Y(n24151) );
  INVXL U17663 ( .A(n24151), .Y(n33863) );
  NOR2X1 U17664 ( .A(n22827), .B(n22825), .Y(n29311) );
  INVXL U17665 ( .A(n24288), .Y(n34325) );
  NOR2BXL U17666 ( .AN(n35422), .B(n35423), .Y(n27965) );
  OAI2BB1XL U17667 ( .A0N(n29257), .A1N(n29676), .B0(n24673), .Y(n27966) );
  INVXL U17668 ( .A(n29364), .Y(n29339) );
  INVXL U17669 ( .A(n27966), .Y(n35426) );
  ADDFXL U17670 ( .A(conv_1[265]), .B(n30191), .CI(n30190), .CO(n29350), .S(
        n30192) );
  AOI2BB1XL U17671 ( .A0N(conv_1[264]), .A1N(n29228), .B0(n29227), .Y(n30190)
         );
  AOI2BB1XL U17672 ( .A0N(conv_1[263]), .A1N(n29280), .B0(n29229), .Y(n29228)
         );
  AOI2BB1XL U17673 ( .A0N(conv_1[261]), .A1N(n29202), .B0(n29229), .Y(n27564)
         );
  INVXL U17674 ( .A(n30191), .Y(n29229) );
  AOI2BB1XL U17675 ( .A0N(conv_1[260]), .A1N(n27560), .B0(n29229), .Y(n29202)
         );
  NOR2X1 U17676 ( .A(n27562), .B(n27561), .Y(n29203) );
  AND2XL U17677 ( .A(n30191), .B(n24693), .Y(n27560) );
  NOR2X1 U17678 ( .A(n30191), .B(n24693), .Y(n27562) );
  AOI21XL U17679 ( .A0(n29233), .A1(n29676), .B0(n18856), .Y(n34080) );
  AOI2BB1XL U17680 ( .A0N(conv_1[250]), .A1N(n35412), .B0(n35414), .Y(n26970)
         );
  AOI2BB1XL U17681 ( .A0N(conv_1[249]), .A1N(n35411), .B0(n35414), .Y(n35412)
         );
  INVXL U17682 ( .A(n33663), .Y(n35414) );
  OAI2BB1XL U17683 ( .A0N(n27987), .A1N(n29676), .B0(n24673), .Y(n33658) );
  NOR2X1 U17684 ( .A(n33423), .B(n33536), .Y(n33533) );
  INVXL U17685 ( .A(n33658), .Y(n35417) );
  OAI2BB1XL U17686 ( .A0N(n33852), .A1N(n29676), .B0(n24208), .Y(n23362) );
  INVXL U17687 ( .A(n23362), .Y(n35408) );
  AOI2BB1XL U17688 ( .A0N(conv_1[220]), .A1N(n25437), .B0(n28602), .Y(n28599)
         );
  INVXL U17689 ( .A(n35392), .Y(n28602) );
  INVXL U17690 ( .A(n24293), .Y(n35395) );
  NOR2BXL U17691 ( .AN(n35385), .B(conv_1[206]), .Y(n35387) );
  NAND2XL U17692 ( .A(n27632), .B(n27849), .Y(n34060) );
  NOR2X1 U17693 ( .A(n23444), .B(n23443), .Y(n23682) );
  INVXL U17694 ( .A(n34060), .Y(n35379) );
  AOI2BB1XL U17695 ( .A0N(conv_1[200]), .A1N(n23445), .B0(n34060), .Y(n23680)
         );
  OAI2BB1XL U17696 ( .A0N(n33122), .A1N(n29676), .B0(n24673), .Y(n35374) );
  AND2XL U17697 ( .A(n35379), .B(n23439), .Y(n23445) );
  INVXL U17698 ( .A(n35374), .Y(n35384) );
  AOI2BB1XL U17699 ( .A0N(conv_1[189]), .A1N(n25062), .B0(n32988), .Y(n35363)
         );
  AOI2BB1XL U17700 ( .A0N(conv_1[188]), .A1N(n35357), .B0(n32988), .Y(n25062)
         );
  INVXL U17701 ( .A(n32988), .Y(n35365) );
  AOI21XL U17702 ( .A0(n32995), .A1(n29676), .B0(n18856), .Y(n35368) );
  INVXL U17703 ( .A(n23923), .Y(n27538) );
  NOR2X1 U17704 ( .A(n23923), .B(n27539), .Y(n23922) );
  AOI2BB1XL U17705 ( .A0N(conv_1[156]), .A1N(n23405), .B0(n23406), .Y(n24312)
         );
  OAI2BB1XL U17706 ( .A0N(n23375), .A1N(n29676), .B0(n24673), .Y(n24429) );
  AND2XL U17707 ( .A(n23394), .B(n23298), .Y(n23400) );
  NOR2X1 U17708 ( .A(n23394), .B(n23298), .Y(n23399) );
  INVXL U17709 ( .A(n24429), .Y(n34048) );
  OAI2BB1XL U17710 ( .A0N(n26831), .A1N(n29676), .B0(n24673), .Y(n35341) );
  OAI2BB1XL U17711 ( .A0N(n33047), .A1N(n29676), .B0(n24673), .Y(n23883) );
  INVXL U17712 ( .A(n23883), .Y(n34296) );
  NOR2BXL U17713 ( .AN(n35331), .B(conv_1[116]), .Y(n35333) );
  OAI2BB1XL U17714 ( .A0N(conv_1[115]), .A1N(n34556), .B0(n31344), .Y(n35332)
         );
  INVXL U17715 ( .A(n34557), .Y(n31344) );
  ADDFXL U17716 ( .A(conv_1[112]), .B(n34557), .CI(n25091), .CO(n31343), .S(
        n24350) );
  AOI2BB1XL U17717 ( .A0N(conv_1[111]), .A1N(n31349), .B0(n31350), .Y(n25091)
         );
  OAI2BB1XL U17718 ( .A0N(n29261), .A1N(n29676), .B0(n24673), .Y(n25090) );
  AOI2BB1XL U17719 ( .A0N(conv_1[110]), .A1N(n29292), .B0(n31344), .Y(n31349)
         );
  AOI2BB1XL U17720 ( .A0N(n29297), .A1N(n29293), .B0(n34557), .Y(n31350) );
  NOR2X1 U17721 ( .A(n31344), .B(n24349), .Y(n29292) );
  AND2XL U17722 ( .A(n31344), .B(n24349), .Y(n29293) );
  AOI22XL U17723 ( .A0(n35181), .A1(n22844), .B0(n28414), .B1(n22843), .Y(
        n22854) );
  AOI22XL U17724 ( .A0(n35130), .A1(n22849), .B0(n34827), .B1(n22848), .Y(
        n22852) );
  INVXL U17725 ( .A(n25090), .Y(n35330) );
  INVXL U17726 ( .A(n31334), .Y(n31337) );
  NAND2XL U17727 ( .A(n27632), .B(n34450), .Y(n31334) );
  AND2XL U17728 ( .A(n31337), .B(n26514), .Y(n26779) );
  NOR2X1 U17729 ( .A(n31337), .B(n26514), .Y(n26778) );
  INVXL U17730 ( .A(n26515), .Y(n31361) );
  OAI2BB1XL U17731 ( .A0N(n26838), .A1N(n29676), .B0(n24673), .Y(n24342) );
  NOR2X1 U17732 ( .A(n22869), .B(n22871), .Y(n34052) );
  INVXL U17733 ( .A(n24342), .Y(n34057) );
  NOR2X1 U17734 ( .A(n27099), .B(n27095), .Y(n33637) );
  AOI2BB1XL U17735 ( .A0N(conv_1[69]), .A1N(n27094), .B0(n35324), .Y(n33635)
         );
  NOR2X1 U17736 ( .A(n27200), .B(n35324), .Y(n27094) );
  NOR2X1 U17737 ( .A(conv_1[68]), .B(n27199), .Y(n27200) );
  NOR2X1 U17738 ( .A(n35326), .B(n35323), .Y(n27201) );
  AOI2BB1XL U17739 ( .A0N(conv_1[67]), .A1N(n35322), .B0(n35324), .Y(n27199)
         );
  OAI2BB1XL U17740 ( .A0N(n27211), .A1N(n29676), .B0(n24673), .Y(n33633) );
  NAND2XL U17741 ( .A(n27632), .B(n34699), .Y(n35324) );
  AOI2BB1XL U17742 ( .A0N(conv_1[66]), .A1N(n27100), .B0(n35324), .Y(n35322)
         );
  NOR2X1 U17743 ( .A(n35324), .B(n26141), .Y(n27107) );
  AND2XL U17744 ( .A(n35324), .B(n26141), .Y(n27106) );
  INVXL U17745 ( .A(n33633), .Y(n35327) );
  NOR2X1 U17746 ( .A(n26824), .B(n27312), .Y(n27317) );
  AOI21XL U17747 ( .A0(n33054), .A1(n29676), .B0(n18856), .Y(n35319) );
  OAI2BB1XL U17748 ( .A0N(n33127), .A1N(n29676), .B0(n24673), .Y(n25080) );
  AOI2BB1XL U17749 ( .A0N(conv_1[39]), .A1N(n27306), .B0(n35289), .Y(n35294)
         );
  AND2XL U17750 ( .A(n35296), .B(n25079), .Y(n27294) );
  NOR2X1 U17751 ( .A(n35296), .B(n25079), .Y(n27295) );
  INVXL U17752 ( .A(n25080), .Y(n35302) );
  INVXL U17753 ( .A(n35296), .Y(n35289) );
  AOI2BB1XL U17754 ( .A0N(conv_1[25]), .A1N(n35273), .B0(n30588), .Y(n30586)
         );
  NOR2X1 U17755 ( .A(n27611), .B(n27610), .Y(n35274) );
  NAND2XL U17756 ( .A(n34721), .B(n27632), .Y(n30588) );
  INVXL U17757 ( .A(n30588), .Y(n35275) );
  AND2XL U17758 ( .A(n35275), .B(n26505), .Y(n27332) );
  AOI21XL U17759 ( .A0(n33443), .A1(n29676), .B0(n18856), .Y(n35278) );
  NOR2X1 U17760 ( .A(conv_1[11]), .B(n26298), .Y(n24538) );
  NOR2X1 U17761 ( .A(n24542), .B(n24540), .Y(n26297) );
  INVXL U17762 ( .A(n24536), .Y(n34552) );
  OR4XL U17763 ( .A(n26298), .B(n34547), .C(conv_1[11]), .D(conv_1[12]), .Y(
        n27363) );
  NOR2X1 U17764 ( .A(conv_2[535]), .B(n33371), .Y(n33372) );
  NOR2X1 U17765 ( .A(n29099), .B(n29094), .Y(n33373) );
  AOI2BB1XL U17766 ( .A0N(conv_2[534]), .A1N(n29093), .B0(n29095), .Y(n33371)
         );
  NOR2X1 U17767 ( .A(n33627), .B(n29095), .Y(n29093) );
  AOI2BB1XL U17768 ( .A0N(conv_2[529]), .A1N(n28852), .B0(n28853), .Y(n30982)
         );
  OAI2BB1XL U17769 ( .A0N(n30427), .A1N(n29676), .B0(n24673), .Y(n33624) );
  OAI21XL U17770 ( .A0(n35229), .A1(n26112), .B0(n35227), .Y(n34926) );
  AOI222XL U17771 ( .A0(n26111), .A1(n26110), .B0(n26111), .B1(n26109), .C0(
        n26110), .C1(n26108), .Y(n26112) );
  AOI22XL U17772 ( .A0(n36245), .A1(n25459), .B0(n25464), .B1(n26374), .Y(
        n34927) );
  OAI21XL U17773 ( .A0(n35229), .A1(n18450), .B0(n35227), .Y(n34940) );
  AOI222XL U17774 ( .A0(n18449), .A1(n18448), .B0(n18449), .B1(n18447), .C0(
        n18448), .C1(n18446), .Y(n18450) );
  INVXL U17775 ( .A(n33624), .Y(n34496) );
  NAND2XL U17776 ( .A(n33580), .B(n27770), .Y(n28202) );
  NOR2X1 U17777 ( .A(n28704), .B(n28706), .Y(n27793) );
  NOR2X1 U17778 ( .A(n28708), .B(n28707), .Y(n27794) );
  AOI2BB1XL U17779 ( .A0N(conv_2[518]), .A1N(n27781), .B0(n28706), .Y(n28705)
         );
  INVXL U17780 ( .A(n28706), .Y(n33580) );
  OAI2BB1XL U17781 ( .A0N(n29443), .A1N(n29676), .B0(n24673), .Y(n33575) );
  INVXL U17782 ( .A(n33575), .Y(n31013) );
  INVXL U17783 ( .A(n36081), .Y(n36088) );
  AOI21XL U17784 ( .A0(n34016), .A1(n29676), .B0(n18856), .Y(n36091) );
  AOI2BB1XL U17785 ( .A0N(conv_2[487]), .A1N(n27758), .B0(n27759), .Y(n30863)
         );
  OAI2BB1XL U17786 ( .A0N(n34670), .A1N(n29676), .B0(n24673), .Y(n33598) );
  AND2XL U17787 ( .A(n34132), .B(n27741), .Y(n27745) );
  INVXL U17788 ( .A(n33598), .Y(n34137) );
  AOI2BB1XL U17789 ( .A0N(conv_2[473]), .A1N(n27879), .B0(n27943), .Y(n30901)
         );
  AOI21XL U17790 ( .A0(n33896), .A1(n33892), .B0(n27943), .Y(n27872) );
  AOI21XL U17791 ( .A0(n27950), .A1(n29676), .B0(n18856), .Y(n34177) );
  NOR2X1 U17792 ( .A(n33609), .B(n27677), .Y(n27660) );
  NOR2X1 U17793 ( .A(conv_2[460]), .B(n33608), .Y(n33609) );
  NOR2X1 U17794 ( .A(n27655), .B(n27654), .Y(n33610) );
  OAI2BB1XL U17795 ( .A0N(n27964), .A1N(n29676), .B0(n24208), .Y(n33606) );
  ADDFXL U17796 ( .A(conv_2[454]), .B(n27643), .CI(n27642), .CO(n30876), .S(
        n24339) );
  INVXL U17797 ( .A(n33606), .Y(n34441) );
  INVXL U17798 ( .A(n28937), .Y(n36067) );
  NAND2XL U17799 ( .A(n34224), .B(n28739), .Y(n28937) );
  AND2XL U17800 ( .A(n36067), .B(n27905), .Y(n28943) );
  NOR2X1 U17801 ( .A(n36067), .B(n27905), .Y(n28942) );
  AOI21XL U17802 ( .A0(n27927), .A1(n29676), .B0(n18856), .Y(n36070) );
  ADDFXL U17803 ( .A(conv_2[430]), .B(n34211), .CI(n32891), .CO(n34210), .S(
        n32892) );
  NOR2BXL U17804 ( .AN(n36054), .B(n36055), .Y(n32891) );
  AND2XL U17805 ( .A(n34211), .B(n28133), .Y(n28893) );
  AOI21XL U17806 ( .A0(n28897), .A1(n29676), .B0(n18856), .Y(n36053) );
  ADDFXL U17807 ( .A(conv_2[416]), .B(n36045), .CI(n33320), .CO(n36044), .S(
        n30886) );
  AOI2BB1XL U17808 ( .A0N(n36037), .A1N(conv_2[415]), .B0(n36038), .Y(n33320)
         );
  NOR2X1 U17809 ( .A(n33690), .B(n33321), .Y(n36037) );
  NOR2X1 U17810 ( .A(n30885), .B(n30884), .Y(n33691) );
  AOI2BB1XL U17811 ( .A0N(conv_2[413]), .A1N(n30883), .B0(n33321), .Y(n33689)
         );
  AOI2BB1XL U17812 ( .A0N(conv_2[412]), .A1N(n28082), .B0(n33321), .Y(n30883)
         );
  INVXL U17813 ( .A(n36045), .Y(n33321) );
  OAI2BB1XL U17814 ( .A0N(n33325), .A1N(n29676), .B0(n24208), .Y(n33687) );
  INVXL U17815 ( .A(n33687), .Y(n36047) );
  OAI21XL U17816 ( .A0(n33141), .A1(n33140), .B0(n33953), .Y(n36033) );
  ADDFXL U17817 ( .A(conv_2[397]), .B(n34634), .CI(n29498), .CO(n34635), .S(
        n24452) );
  AOI2BB1XL U17818 ( .A0N(conv_2[396]), .A1N(n28108), .B0(n28109), .Y(n29498)
         );
  OAI2BB1XL U17819 ( .A0N(n33262), .A1N(n29676), .B0(n24208), .Y(n24451) );
  AOI2BB1XL U17820 ( .A0N(conv_2[395]), .A1N(n28114), .B0(n33953), .Y(n28108)
         );
  AOI2BB1XL U17821 ( .A0N(n28119), .A1N(n28115), .B0(n34634), .Y(n28109) );
  INVXL U17822 ( .A(n24451), .Y(n36031) );
  AOI2BB1XL U17823 ( .A0N(conv_2[384]), .A1N(n28012), .B0(n28013), .Y(n28018)
         );
  AOI21XL U17824 ( .A0(n33675), .A1(conv_2[383]), .B0(n34529), .Y(n28013) );
  NOR2X1 U17825 ( .A(n36024), .B(n36027), .Y(n33675) );
  INVXL U17826 ( .A(n34529), .Y(n36025) );
  OAI2BB1XL U17827 ( .A0N(n28160), .A1N(n29676), .B0(n24208), .Y(n34531) );
  AND2XL U17828 ( .A(n34529), .B(n23079), .Y(n29444) );
  INVXL U17829 ( .A(n34531), .Y(n36028) );
  OR4XL U17830 ( .A(n34528), .B(conv_2[387]), .C(conv_2[386]), .D(n36025), .Y(
        n28155) );
  AOI2BB1XL U17831 ( .A0N(conv_2[369]), .A1N(n29492), .B0(n29493), .Y(n27272)
         );
  OAI2BB1XL U17832 ( .A0N(n29472), .A1N(n29676), .B0(n24208), .Y(n24455) );
  OAI211X1 U17833 ( .A0(n22807), .A1(n34989), .B0(n22806), .C0(n22805), .Y(
        n34502) );
  AOI21XL U17834 ( .A0(n28324), .A1(n22802), .B0(n22801), .Y(n22806) );
  AOI22XL U17835 ( .A0(n34827), .A1(n22804), .B0(n16755), .B1(n22803), .Y(
        n22805) );
  OAI2BB2XL U17836 ( .B0(n22800), .B1(n35135), .A0N(n23240), .A1N(n16670), .Y(
        n22801) );
  INVXL U17837 ( .A(n24455), .Y(n36017) );
  INVXL U17838 ( .A(n29526), .Y(n33925) );
  OAI31XL U17839 ( .A0(conv_2[352]), .A1(conv_2[353]), .A2(n29523), .B0(n29526), .Y(n27995) );
  NOR2X1 U17840 ( .A(n29526), .B(n29523), .Y(n29518) );
  OAI2BB1XL U17841 ( .A0N(n29465), .A1N(n29676), .B0(n24208), .Y(n24190) );
  AOI22XL U17842 ( .A0(n26470), .A1(n23092), .B0(n34827), .B1(n23091), .Y(
        n23093) );
  AOI22XL U17843 ( .A0(n28465), .A1(n23090), .B0(n16755), .B1(n23089), .Y(
        n23094) );
  INVXL U17844 ( .A(n24190), .Y(n36010) );
  INVXL U17845 ( .A(n35995), .Y(n35997) );
  NOR2X1 U17846 ( .A(n35995), .B(n35996), .Y(n28103) );
  OAI2BB1XL U17847 ( .A0N(n29453), .A1N(n29676), .B0(n24208), .Y(n24303) );
  OAI2BB1XL U17848 ( .A0N(n33237), .A1N(n29676), .B0(n24208), .Y(n24298) );
  INVXL U17849 ( .A(n24298), .Y(n35986) );
  OAI2BB1XL U17850 ( .A0N(n33985), .A1N(n29676), .B0(n24208), .Y(n34026) );
  AND2XL U17851 ( .A(n33979), .B(n19114), .Y(n30857) );
  INVXL U17852 ( .A(n34026), .Y(n35976) );
  AOI2BB1XL U17853 ( .A0N(conv_2[292]), .A1N(n30917), .B0(n30916), .Y(n30999)
         );
  OAI2BB1XL U17854 ( .A0N(n33300), .A1N(n29676), .B0(n24208), .Y(n35959) );
  AND2XL U17855 ( .A(n35957), .B(n28091), .Y(n30888) );
  INVXL U17856 ( .A(n35959), .Y(n35963) );
  NOR2X1 U17857 ( .A(n28883), .B(n18955), .Y(n28007) );
  OAI2BB1XL U17858 ( .A0N(n28890), .A1N(n29676), .B0(n24208), .Y(n35952) );
  AOI2BB1XL U17859 ( .A0N(conv_2[260]), .A1N(n28177), .B0(n28161), .Y(n34599)
         );
  AOI2BB1XL U17860 ( .A0N(n28182), .A1N(n28178), .B0(n28191), .Y(n34600) );
  NOR2X1 U17861 ( .A(n28161), .B(n19043), .Y(n28177) );
  AOI21XL U17862 ( .A0(n28144), .A1(n29676), .B0(n18856), .Y(n34601) );
  AOI22XL U17863 ( .A0(n34827), .A1(n23089), .B0(n16755), .B1(n22403), .Y(
        n19037) );
  NOR2X1 U17864 ( .A(conv_2[249]), .B(n33681), .Y(n33682) );
  NOR2X1 U17865 ( .A(n29154), .B(n29150), .Y(n33683) );
  AOI2BB1XL U17866 ( .A0N(conv_2[248]), .A1N(n29149), .B0(n29455), .Y(n33681)
         );
  OAI2BB1XL U17867 ( .A0N(n28153), .A1N(n29676), .B0(n24208), .Y(n33679) );
  AOI2BB1XL U17868 ( .A0N(conv_2[247]), .A1N(n29167), .B0(n29455), .Y(n29149)
         );
  INVXL U17869 ( .A(n33679), .Y(n35945) );
  OAI2BB1XL U17870 ( .A0N(n33101), .A1N(n29676), .B0(n24208), .Y(n29599) );
  NOR2X1 U17871 ( .A(n32876), .B(n29184), .Y(n29183) );
  AOI2BB1XL U17872 ( .A0N(conv_2[230]), .A1N(n29512), .B0(n33096), .Y(n29173)
         );
  INVXL U17873 ( .A(n29599), .Y(n34458) );
  INVXL U17874 ( .A(n32876), .Y(n33096) );
  NAND2XL U17875 ( .A(conv_2[218]), .B(n33769), .Y(n30428) );
  AOI2BB1XL U17876 ( .A0N(conv_2[217]), .A1N(n30155), .B0(n31121), .Y(n33767)
         );
  NOR2X1 U17877 ( .A(conv_2[218]), .B(n33767), .Y(n33768) );
  NOR2X1 U17878 ( .A(n30154), .B(n30159), .Y(n33769) );
  NOR2X1 U17879 ( .A(n33770), .B(n30155), .Y(n30154) );
  OAI2BB1XL U17880 ( .A0N(n31126), .A1N(n29676), .B0(n24208), .Y(n33765) );
  OAI2BB1XL U17881 ( .A0N(n33040), .A1N(n29676), .B0(n24208), .Y(n29607) );
  AOI2BB1XL U17882 ( .A0N(conv_2[204]), .A1N(n29927), .B0(n35928), .Y(n29606)
         );
  AOI2BB1XL U17883 ( .A0N(conv_2[203]), .A1N(n35926), .B0(n35928), .Y(n29927)
         );
  INVXL U17884 ( .A(n29935), .Y(n35928) );
  INVXL U17885 ( .A(n29607), .Y(n35931) );
  NOR2X1 U17886 ( .A(n29893), .B(n29892), .Y(n33457) );
  OAI2BB1XL U17887 ( .A0N(n29958), .A1N(n29676), .B0(n24279), .Y(n33453) );
  NOR2X1 U17888 ( .A(n29890), .B(n29886), .Y(n35913) );
  INVXL U17889 ( .A(n30946), .Y(n35914) );
  AND2XL U17890 ( .A(n35914), .B(n28655), .Y(n29898) );
  INVXL U17891 ( .A(n33453), .Y(n35917) );
  OAI2BB1XL U17892 ( .A0N(n34598), .A1N(n29676), .B0(n24279), .Y(n30969) );
  AND2XL U17893 ( .A(n29831), .B(n29834), .Y(n29840) );
  NOR2X1 U17894 ( .A(n29831), .B(n29834), .Y(n29839) );
  INVXL U17895 ( .A(n30969), .Y(n34589) );
  OR3XL U17896 ( .A(n34585), .B(conv_2[177]), .C(n33974), .Y(n34593) );
  OAI31XL U17897 ( .A0(conv_2[157]), .A1(conv_2[158]), .A2(n29863), .B0(n34626), .Y(n34625) );
  OAI2BB1XL U17898 ( .A0N(n24535), .A1N(n29676), .B0(n24279), .Y(n24358) );
  INVXL U17899 ( .A(n35899), .Y(n35907) );
  OAI2BB1XL U17900 ( .A0N(n30239), .A1N(n29676), .B0(n24279), .Y(n35909) );
  AND2XL U17901 ( .A(n35907), .B(n27972), .Y(n34240) );
  NOR2X1 U17902 ( .A(n35907), .B(n27972), .Y(n34239) );
  INVXL U17903 ( .A(n35909), .Y(n35902) );
  AOI2BB1XL U17904 ( .A0N(conv_2[127]), .A1N(n30061), .B0(n30062), .Y(n24361)
         );
  OAI2BB1XL U17905 ( .A0N(n30448), .A1N(n29676), .B0(n24279), .Y(n33801) );
  AND2XL U17906 ( .A(n34344), .B(n24354), .Y(n34124) );
  NOR2X1 U17907 ( .A(n34344), .B(n24354), .Y(n34125) );
  INVXL U17908 ( .A(n33801), .Y(n34491) );
  INVXL U17909 ( .A(n34344), .Y(n30443) );
  AOI2BB1XL U17910 ( .A0N(conv_2[113]), .A1N(n35889), .B0(n35884), .Y(n28682)
         );
  AOI2BB1XL U17911 ( .A0N(conv_2[112]), .A1N(n35882), .B0(n35884), .Y(n35889)
         );
  NOR2X1 U17912 ( .A(n35886), .B(n35883), .Y(n35890) );
  NAND2XL U17913 ( .A(n28739), .B(n34717), .Y(n35884) );
  INVXL U17914 ( .A(n23575), .Y(n35894) );
  NOR2X1 U17915 ( .A(n30218), .B(n30216), .Y(n30226) );
  INVXL U17916 ( .A(n23033), .Y(n34447) );
  NOR2X1 U17917 ( .A(conv_2[86]), .B(n31003), .Y(n30927) );
  NOR2X1 U17918 ( .A(conv_2[85]), .B(n33811), .Y(n33812) );
  NOR2X1 U17919 ( .A(n30174), .B(n30173), .Y(n33813) );
  OAI2BB1XL U17920 ( .A0N(n32677), .A1N(n29676), .B0(n24279), .Y(n33809) );
  NOR2X1 U17921 ( .A(conv_2[84]), .B(n28744), .Y(n30172) );
  NOR2X1 U17922 ( .A(n30171), .B(n30167), .Y(n35875) );
  NAND2XL U17923 ( .A(n28739), .B(n34438), .Y(n30924) );
  INVXL U17924 ( .A(n30924), .Y(n35876) );
  AND2XL U17925 ( .A(n35876), .B(n28742), .Y(n30179) );
  NOR2X1 U17926 ( .A(n35876), .B(n28742), .Y(n30178) );
  INVXL U17927 ( .A(n33809), .Y(n35879) );
  NOR2X1 U17928 ( .A(n30243), .B(n30241), .Y(n33734) );
  AND2XL U17929 ( .A(n33735), .B(n30106), .Y(n30118) );
  NAND2BXL U17930 ( .AN(conv_2[67]), .B(n18972), .Y(n30106) );
  OAI21XL U17931 ( .A0(conv_2[66]), .A1(n30100), .B0(n33735), .Y(n18972) );
  NOR2X1 U17932 ( .A(n30105), .B(n30101), .Y(n30107) );
  NOR2XL U17933 ( .A(n29830), .B(n31418), .Y(n33735) );
  OAI2BB1XL U17934 ( .A0N(n30247), .A1N(n29676), .B0(n24279), .Y(n33730) );
  AOI2BB1XL U17935 ( .A0N(conv_2[65]), .A1N(n30112), .B0(n30242), .Y(n30100)
         );
  INVXL U17936 ( .A(n33735), .Y(n30242) );
  INVXL U17937 ( .A(n33730), .Y(n35846) );
  AOI2BB1XL U17938 ( .A0N(conv_2[53]), .A1N(n27814), .B0(n31134), .Y(n28713)
         );
  INVXL U17939 ( .A(n31137), .Y(n31134) );
  OAI2BB1XL U17940 ( .A0N(n33108), .A1N(n29676), .B0(n24279), .Y(n30873) );
  AOI2BB1XL U17941 ( .A0N(conv_2[50]), .A1N(n27806), .B0(n31134), .Y(n27819)
         );
  INVXL U17942 ( .A(n30873), .Y(n34505) );
  NOR2X1 U17943 ( .A(n35864), .B(n35861), .Y(n33587) );
  AOI2BB1XL U17944 ( .A0N(conv_2[39]), .A1N(n35860), .B0(n35862), .Y(n33585)
         );
  AOI2BB1XL U17945 ( .A0N(conv_2[38]), .A1N(n27717), .B0(n35862), .Y(n35860)
         );
  INVXL U17946 ( .A(n35862), .Y(n33588) );
  INVXL U17947 ( .A(n33986), .Y(n35865) );
  OAI2BB1XL U17948 ( .A0N(n27957), .A1N(n29676), .B0(n24279), .Y(n33986) );
  NOR2X1 U17949 ( .A(n27916), .B(n28673), .Y(n27837) );
  NOR2X1 U17950 ( .A(conv_2[25]), .B(n27915), .Y(n27916) );
  NOR2X1 U17951 ( .A(n28675), .B(n28674), .Y(n27917) );
  NOR2X1 U17952 ( .A(n28671), .B(n28673), .Y(n27915) );
  NOR2X1 U17953 ( .A(n33618), .B(n28673), .Y(n28672) );
  NOR2X1 U17954 ( .A(conv_2[24]), .B(n28672), .Y(n28671) );
  NOR2X1 U17955 ( .A(conv_2[23]), .B(n33617), .Y(n33618) );
  NOR2X1 U17956 ( .A(n27830), .B(n28673), .Y(n33617) );
  OAI2BB1XL U17957 ( .A0N(n27942), .A1N(n29676), .B0(n24279), .Y(n33615) );
  AOI2BB1XL U17958 ( .A0N(conv_2[21]), .A1N(n29082), .B0(n28673), .Y(n27557)
         );
  NOR2X1 U17959 ( .A(conv_2[22]), .B(n27557), .Y(n27830) );
  INVXL U17960 ( .A(n33615), .Y(n30412) );
  OAI2BB1XL U17961 ( .A0N(n27935), .A1N(n29676), .B0(n24279), .Y(n33566) );
  INVXL U17962 ( .A(n33566), .Y(n30958) );
  NOR2X1 U17963 ( .A(conv_3[534]), .B(n28958), .Y(n28957) );
  NOR2X1 U17964 ( .A(conv_3[533]), .B(n33716), .Y(n33717) );
  NOR2X1 U17965 ( .A(n27571), .B(n27570), .Y(n33718) );
  INVXL U17966 ( .A(n33719), .Y(n28959) );
  NOR2X1 U17967 ( .A(conv_3[532]), .B(n27569), .Y(n27568) );
  AOI2BB1XL U17968 ( .A0N(conv_3[529]), .A1N(n24365), .B0(n24364), .Y(n26302)
         );
  OAI2BB1XL U17969 ( .A0N(n31290), .A1N(n29676), .B0(n25246), .Y(n33714) );
  INVXL U17970 ( .A(n23783), .Y(n34969) );
  AOI22XL U17971 ( .A0(n34963), .A1(n34962), .B0(n34961), .B1(n34960), .Y(
        n34967) );
  OAI21XL U17972 ( .A0(n35229), .A1(n20596), .B0(n35227), .Y(n34978) );
  AOI222XL U17973 ( .A0(n20595), .A1(n20594), .B0(n20595), .B1(n20593), .C0(
        n20594), .C1(n20592), .Y(n20596) );
  INVXL U17974 ( .A(n26451), .Y(n34983) );
  OAI2BB1XL U17975 ( .A0N(n28391), .A1N(n24903), .B0(n35227), .Y(n35001) );
  AOI222XL U17976 ( .A0(n24902), .A1(n24901), .B0(n24902), .B1(n24900), .C0(
        n24901), .C1(n24899), .Y(n24903) );
  AOI211XL U17977 ( .A0(n26470), .A1(n35175), .B0(n24818), .C0(n24817), .Y(
        n24902) );
  AOI211XL U17978 ( .A0(n22762), .A1(conv_3[75]), .B0(n22243), .C0(n22242), 
        .Y(n35240) );
  NOR2X1 U17979 ( .A(n24039), .B(n30832), .Y(n22243) );
  OAI21XL U17980 ( .A0(n35229), .A1(n35228), .B0(n35227), .Y(n35250) );
  INVXL U17981 ( .A(n33714), .Y(n31191) );
  ADDFXL U17982 ( .A(conv_3[520]), .B(n31180), .CI(n26677), .CO(n31292), .S(
        n24480) );
  AOI2BB1XL U17983 ( .A0N(conv_3[519]), .A1N(n31147), .B0(n31148), .Y(n26677)
         );
  AOI21XL U17984 ( .A0(n31179), .A1(conv_3[518]), .B0(n31180), .Y(n31148) );
  OAI2BB1XL U17985 ( .A0N(n31296), .A1N(n29676), .B0(n29675), .Y(n24479) );
  OAI211X1 U17986 ( .A0(n23252), .A1(n34989), .B0(n23251), .C0(n23250), .Y(
        n34019) );
  AOI21XL U17987 ( .A0(n34827), .A1(n23249), .B0(n23248), .Y(n23250) );
  OAI211XL U17988 ( .A0(n23247), .A1(n35159), .B0(n23246), .C0(n23245), .Y(
        n23248) );
  INVXL U17989 ( .A(n24479), .Y(n33303) );
  OR4XL U17990 ( .A(n31292), .B(conv_3[521]), .C(conv_3[522]), .D(n31291), .Y(
        n33301) );
  INVXL U17991 ( .A(n33918), .Y(n35838) );
  AND2XL U17992 ( .A(n35838), .B(n27627), .Y(n32071) );
  NOR2X1 U17993 ( .A(n35838), .B(n27627), .Y(n32070) );
  AOI21XL U17994 ( .A0(n34519), .A1(n29676), .B0(n18856), .Y(n35841) );
  OR2XL U17995 ( .A(n35831), .B(n35822), .Y(n35817) );
  OAI2BB1XL U17996 ( .A0N(n32233), .A1N(n29676), .B0(n29675), .Y(n35833) );
  AOI21XL U17997 ( .A0(n23055), .A1(n23273), .B0(n23054), .Y(n23056) );
  INVXL U17998 ( .A(n35833), .Y(n35826) );
  INVXL U17999 ( .A(n35810), .Y(n32328) );
  AOI2BB1XL U18000 ( .A0N(conv_3[475]), .A1N(n32185), .B0(n32328), .Y(n32339)
         );
  OAI2BB1XL U18001 ( .A0N(conv_3[475]), .A1N(n32185), .B0(n32328), .Y(n32340)
         );
  AOI2BB1XL U18002 ( .A0N(conv_3[471]), .A1N(n35808), .B0(n32328), .Y(n32333)
         );
  AOI21XL U18003 ( .A0(n35809), .A1(conv_3[471]), .B0(n35810), .Y(n32334) );
  AOI2BB1XL U18004 ( .A0N(conv_3[470]), .A1N(n26120), .B0(n32328), .Y(n35808)
         );
  NOR2X1 U18005 ( .A(n26121), .B(n26124), .Y(n35809) );
  AND2XL U18006 ( .A(n35810), .B(n19021), .Y(n26120) );
  AOI21XL U18007 ( .A0(n32189), .A1(n29676), .B0(n18856), .Y(n35813) );
  AOI2BB1XL U18008 ( .A0N(conv_3[460]), .A1N(n31513), .B0(n31517), .Y(n31523)
         );
  ADDFXL U18009 ( .A(conv_3[459]), .B(n33780), .CI(n32594), .CO(n31513), .S(
        n32595) );
  AOI2BB1XL U18010 ( .A0N(n35801), .A1N(conv_3[458]), .B0(n35802), .Y(n32594)
         );
  NOR2X1 U18011 ( .A(n33777), .B(n31517), .Y(n35801) );
  AOI21XL U18012 ( .A0(n33779), .A1(conv_3[457]), .B0(n33780), .Y(n35802) );
  NOR2X1 U18013 ( .A(n31508), .B(n31512), .Y(n33779) );
  OAI2BB1XL U18014 ( .A0N(n32247), .A1N(n29676), .B0(n29675), .Y(n33774) );
  AOI2BB1XL U18015 ( .A0N(conv_3[456]), .A1N(n31507), .B0(n31517), .Y(n33776)
         );
  NOR2X1 U18016 ( .A(n35798), .B(n31517), .Y(n31507) );
  NOR2X1 U18017 ( .A(conv_3[445]), .B(n33758), .Y(n33759) );
  NOR2X1 U18018 ( .A(n35791), .B(n35788), .Y(n33760) );
  AOI2BB1XL U18019 ( .A0N(conv_3[444]), .A1N(n35787), .B0(n35789), .Y(n33758)
         );
  NOR2X1 U18020 ( .A(n32109), .B(n35789), .Y(n35787) );
  NOR2X1 U18021 ( .A(conv_3[443]), .B(n32108), .Y(n32109) );
  NOR2X1 U18022 ( .A(n35784), .B(n35782), .Y(n32110) );
  INVXL U18023 ( .A(n35789), .Y(n33761) );
  AOI2BB1XL U18024 ( .A0N(conv_3[442]), .A1N(n35781), .B0(n35789), .Y(n32108)
         );
  OAI2BB1XL U18025 ( .A0N(n32149), .A1N(n29676), .B0(n29675), .Y(n33756) );
  AOI2BB1XL U18026 ( .A0N(conv_3[441]), .A1N(n31938), .B0(n35789), .Y(n35781)
         );
  NAND2XL U18027 ( .A(n31924), .B(n34224), .Y(n35789) );
  AND2XL U18028 ( .A(n33761), .B(n31927), .Y(n31933) );
  NOR2X1 U18029 ( .A(n33761), .B(n31927), .Y(n31932) );
  INVXL U18030 ( .A(n33756), .Y(n35792) );
  AOI2BB1XL U18031 ( .A0N(conv_3[430]), .A1N(n31726), .B0(n35775), .Y(n32157)
         );
  NAND2XL U18032 ( .A(n31924), .B(n34768), .Y(n35775) );
  OAI2BB1XL U18033 ( .A0N(n32162), .A1N(n29676), .B0(n29675), .Y(n33784) );
  INVXL U18034 ( .A(n35775), .Y(n33790) );
  AND2XL U18035 ( .A(n33790), .B(n31696), .Y(n32576) );
  NOR2X1 U18036 ( .A(n33790), .B(n31696), .Y(n32575) );
  INVXL U18037 ( .A(n33784), .Y(n35778) );
  AOI2BB1XL U18038 ( .A0N(conv_3[415]), .A1N(n31993), .B0(n32558), .Y(n32011)
         );
  OAI21XL U18039 ( .A0(n31987), .A1(n31992), .B0(n31988), .Y(n32545) );
  OAI2BB1XL U18040 ( .A0N(n32196), .A1N(n29676), .B0(n29675), .Y(n32546) );
  NOR2X1 U18041 ( .A(n32558), .B(n19206), .Y(n32627) );
  AOI2BB1XL U18042 ( .A0N(conv_3[400]), .A1N(n32050), .B0(n33695), .Y(n33220)
         );
  AOI2BB1XL U18043 ( .A0N(conv_3[397]), .A1N(n32038), .B0(n32037), .Y(n32531)
         );
  OAI2BB1XL U18044 ( .A0N(n34009), .A1N(n29676), .B0(n29675), .Y(n32532) );
  AND2XL U18045 ( .A(n33699), .B(n32020), .Y(n32026) );
  NOR2X1 U18046 ( .A(n33699), .B(n32020), .Y(n32025) );
  INVXL U18047 ( .A(n32532), .Y(n33703) );
  ADDFHX1 U18048 ( .A(conv_3[381]), .B(n34164), .CI(n32622), .CO(n19194), .S(
        n32624) );
  AOI21XL U18049 ( .A0(n31459), .A1(n19193), .B0(n31454), .Y(n32622) );
  NAND2XL U18050 ( .A(n34164), .B(n31455), .Y(n19193) );
  OAI2BB1XL U18051 ( .A0N(n32204), .A1N(n29676), .B0(n29675), .Y(n32623) );
  INVXL U18052 ( .A(n32623), .Y(n34168) );
  INVXL U18053 ( .A(n27532), .Y(n27535) );
  NAND3XL U18054 ( .A(n34164), .B(n34169), .C(n34162), .Y(n34138) );
  NOR2X1 U18055 ( .A(n33831), .B(n35761), .Y(n31631) );
  NOR2X1 U18056 ( .A(n35763), .B(n35760), .Y(n33832) );
  INVXL U18057 ( .A(n35761), .Y(n33833) );
  AOI2BB1XL U18058 ( .A0N(conv_3[369]), .A1N(n35759), .B0(n35761), .Y(n33830)
         );
  OAI2BB1XL U18059 ( .A0N(n32127), .A1N(n29676), .B0(n29675), .Y(n33828) );
  AOI2BB1XL U18060 ( .A0N(conv_3[368]), .A1N(n31648), .B0(n35761), .Y(n35759)
         );
  NAND2XL U18061 ( .A(n31924), .B(n34502), .Y(n35761) );
  AND2XL U18062 ( .A(n33833), .B(n31627), .Y(n31637) );
  NOR2X1 U18063 ( .A(n33833), .B(n31627), .Y(n31636) );
  INVXL U18064 ( .A(n33828), .Y(n35764) );
  NOR2X1 U18065 ( .A(n32131), .B(n32129), .Y(n33726) );
  NOR2X1 U18066 ( .A(conv_3[355]), .B(n33472), .Y(n33473) );
  NOR2X1 U18067 ( .A(n31490), .B(n31486), .Y(n33474) );
  AOI2BB1XL U18068 ( .A0N(conv_3[354]), .A1N(n31485), .B0(n32130), .Y(n33472)
         );
  NOR2X1 U18069 ( .A(n33750), .B(n32130), .Y(n31485) );
  OAI2BB1XL U18070 ( .A0N(n32135), .A1N(n29676), .B0(n29675), .Y(n33747) );
  INVXL U18071 ( .A(n33747), .Y(n34746) );
  AOI2BB1XL U18072 ( .A0N(n35753), .A1N(conv_3[336]), .B0(n35754), .Y(n27588)
         );
  AOI21XL U18073 ( .A0(conv_3[335]), .A1(n35749), .B0(n31980), .Y(n35754) );
  OAI2BB1XL U18074 ( .A0N(n32219), .A1N(n29676), .B0(n29675), .Y(n35756) );
  INVXL U18075 ( .A(n35756), .Y(n35748) );
  AOI21XL U18076 ( .A0(n33841), .A1(conv_3[322]), .B0(n33842), .Y(n35740) );
  NOR2X1 U18077 ( .A(n31909), .B(n31908), .Y(n33841) );
  OAI2BB1XL U18078 ( .A0N(n33287), .A1N(n29676), .B0(n29675), .Y(n33837) );
  AOI2BB1XL U18079 ( .A0N(conv_3[320]), .A1N(n31901), .B0(n33281), .Y(n28759)
         );
  NAND2XL U18080 ( .A(conv_3[320]), .B(n31902), .Y(n31909) );
  INVXL U18081 ( .A(n33837), .Y(n35743) );
  OAI2BB1XL U18082 ( .A0N(n33115), .A1N(n29676), .B0(n29675), .Y(n32614) );
  AND2XL U18083 ( .A(n35732), .B(n31406), .Y(n31443) );
  INVXL U18084 ( .A(n32614), .Y(n35736) );
  ADDFXL U18085 ( .A(conv_3[295]), .B(n35720), .CI(n32565), .CO(n34479), .S(
        n32567) );
  NOR2BXL U18086 ( .AN(n35727), .B(n35728), .Y(n32565) );
  OAI2BB1XL U18087 ( .A0N(n32240), .A1N(n29676), .B0(n29675), .Y(n32566) );
  NOR2BXL U18088 ( .AN(n35725), .B(conv_3[294]), .Y(n35728) );
  OAI2BB1XL U18089 ( .A0N(n35719), .A1N(conv_3[293]), .B0(n31896), .Y(n35727)
         );
  NOR2X1 U18090 ( .A(n31883), .B(n31887), .Y(n35719) );
  INVXL U18091 ( .A(n32566), .Y(n35726) );
  OAI2BB1XL U18092 ( .A0N(n32263), .A1N(n29676), .B0(n29675), .Y(n32619) );
  AOI2BB1XL U18093 ( .A0N(conv_3[277]), .A1N(n31750), .B0(n32599), .Y(n31738)
         );
  OAI211X1 U18094 ( .A0(n22807), .A1(n35135), .B0(n18951), .C0(n18950), .Y(
        n34711) );
  INVXL U18095 ( .A(n32619), .Y(n34709) );
  INVXL U18096 ( .A(n33480), .Y(n33478) );
  AOI21XL U18097 ( .A0(n33911), .A1(n29676), .B0(n18856), .Y(n35713) );
  OAI2BB1XL U18098 ( .A0N(n29129), .A1N(n29676), .B0(n29675), .Y(n33545) );
  INVXL U18099 ( .A(n35700), .Y(n35693) );
  AND2XL U18100 ( .A(n35693), .B(n28798), .Y(n34246) );
  INVXL U18101 ( .A(n33545), .Y(n35706) );
  INVXL U18102 ( .A(n33878), .Y(n35673) );
  AND2XL U18103 ( .A(n35673), .B(n26154), .Y(n29162) );
  NOR2X1 U18104 ( .A(n35673), .B(n26154), .Y(n29161) );
  AOI21XL U18105 ( .A0(n33904), .A1(n29676), .B0(n18856), .Y(n35676) );
  NOR2BXL U18106 ( .AN(n35666), .B(conv_3[221]), .Y(n35668) );
  AOI2BB1XL U18107 ( .A0N(conv_3[219]), .A1N(n31536), .B0(n34649), .Y(n31543)
         );
  NOR2X1 U18108 ( .A(n31541), .B(n31537), .Y(n31542) );
  NOR2X1 U18109 ( .A(conv_3[218]), .B(n32057), .Y(n32058) );
  NOR2X1 U18110 ( .A(n31531), .B(n34649), .Y(n32057) );
  AOI2BB1XL U18111 ( .A0N(conv_3[216]), .A1N(n35658), .B0(n34649), .Y(n28833)
         );
  NAND2XL U18112 ( .A(n34476), .B(n31924), .Y(n34649) );
  NOR2X1 U18113 ( .A(conv_3[217]), .B(n28833), .Y(n31531) );
  AOI2BB1XL U18114 ( .A0N(conv_3[215]), .A1N(n28829), .B0(n34649), .Y(n35658)
         );
  NOR2X1 U18115 ( .A(n28831), .B(n28830), .Y(n35659) );
  INVXL U18116 ( .A(n34649), .Y(n35660) );
  OAI2BB1XL U18117 ( .A0N(n32142), .A1N(n29676), .B0(n29675), .Y(n35662) );
  AND2XL U18118 ( .A(n35660), .B(n26526), .Y(n28829) );
  INVXL U18119 ( .A(n35662), .Y(n35665) );
  AOI2BB1XL U18120 ( .A0N(conv_3[203]), .A1N(n34656), .B0(n31848), .Y(n28838)
         );
  INVXL U18121 ( .A(n35653), .Y(n31848) );
  ADDFXL U18122 ( .A(conv_3[202]), .B(n35653), .CI(n28836), .CO(n34656), .S(
        n24476) );
  AOI2BB1XL U18123 ( .A0N(conv_3[201]), .A1N(n31865), .B0(n31866), .Y(n28836)
         );
  OAI2BB1XL U18124 ( .A0N(n32277), .A1N(n29676), .B0(n22138), .Y(n35655) );
  NOR2X1 U18125 ( .A(n31848), .B(n24475), .Y(n35644) );
  NOR2X1 U18126 ( .A(conv_3[200]), .B(n35644), .Y(n35648) );
  INVXL U18127 ( .A(n35655), .Y(n35646) );
  OAI2BB1XL U18128 ( .A0N(n32212), .A1N(n29676), .B0(n22138), .Y(n32650) );
  AND2XL U18129 ( .A(n32649), .B(n26317), .Y(n31614) );
  AOI22XL U18130 ( .A0(n28414), .A1(n22170), .B0(n35181), .B1(n22122), .Y(
        n22126) );
  INVXL U18131 ( .A(n32650), .Y(n34704) );
  AOI2BB1XL U18132 ( .A0N(conv_3[191]), .A1N(n31621), .B0(n31620), .Y(n32632)
         );
  AOI2BB1XL U18133 ( .A0N(conv_3[170]), .A1N(n31584), .B0(n32221), .Y(n31568)
         );
  NOR2X1 U18134 ( .A(n31585), .B(n31589), .Y(n31567) );
  AND2XL U18135 ( .A(n35639), .B(n31562), .Y(n31584) );
  INVXL U18136 ( .A(n32252), .Y(n32316) );
  AND2XL U18137 ( .A(n32316), .B(n29747), .Y(n32285) );
  AOI21XL U18138 ( .A0(n32256), .A1(n29676), .B0(n18856), .Y(n34751) );
  NOR2X1 U18139 ( .A(n31712), .B(n31708), .Y(n33465) );
  AOI2BB1XL U18140 ( .A0N(conv_3[144]), .A1N(n31707), .B0(n32789), .Y(n33463)
         );
  AOI2BB1XL U18141 ( .A0N(conv_3[143]), .A1N(n31720), .B0(n32789), .Y(n31707)
         );
  INVXL U18142 ( .A(n33466), .Y(n32789) );
  NOR2X1 U18143 ( .A(n33466), .B(n31720), .Y(n31719) );
  OAI2BB1XL U18144 ( .A0N(n32175), .A1N(n29676), .B0(n25246), .Y(n33461) );
  AOI21XL U18145 ( .A0(n34400), .A1(n34395), .B0(n32789), .Y(n31713) );
  OAI211X1 U18146 ( .A0(n19124), .A1(n26409), .B0(n19123), .C0(n19122), .Y(
        n34740) );
  AOI22XL U18147 ( .A0(N18471), .A1(n22267), .B0(n34906), .B1(n22153), .Y(
        n19122) );
  INVXL U18148 ( .A(n33461), .Y(n34737) );
  AOI2BB1XL U18149 ( .A0N(conv_3[128]), .A1N(n31412), .B0(n34783), .Y(n28953)
         );
  OAI2BB1XL U18150 ( .A0N(n34788), .A1N(n29676), .B0(n25246), .Y(n35572) );
  AND2XL U18151 ( .A(n35622), .B(n28951), .Y(n31398) );
  INVXL U18152 ( .A(n35572), .Y(n35626) );
  AOI2BB1XL U18153 ( .A0N(conv_3[131]), .A1N(n33710), .B0(n33709), .Y(n34757)
         );
  INVXL U18154 ( .A(n35622), .Y(n34783) );
  AOI2BB1XL U18155 ( .A0N(conv_3[113]), .A1N(n31791), .B0(n31792), .Y(n32653)
         );
  OAI2BB1XL U18156 ( .A0N(n32270), .A1N(n29676), .B0(n25246), .Y(n32654) );
  INVXL U18157 ( .A(n32654), .Y(n34200) );
  AOI2BB1XL U18158 ( .A0N(conv_3[99]), .A1N(n35613), .B0(n35615), .Y(n32115)
         );
  AOI2BB1XL U18159 ( .A0N(conv_3[98]), .A1N(n31685), .B0(n35615), .Y(n35613)
         );
  NAND2XL U18160 ( .A(n34450), .B(n31924), .Y(n35615) );
  INVXL U18161 ( .A(n16658), .Y(n33912) );
  OAI2BB1XL U18162 ( .A0N(n32120), .A1N(n29676), .B0(n25246), .Y(n33739) );
  INVXL U18163 ( .A(n35615), .Y(n34186) );
  INVXL U18164 ( .A(n33739), .Y(n35618) );
  INVXL U18165 ( .A(n35607), .Y(n31842) );
  AND2XL U18166 ( .A(n31842), .B(n31805), .Y(n34151) );
  NOR2X1 U18167 ( .A(n31842), .B(n31805), .Y(n34150) );
  NAND4X1 U18168 ( .A(n22407), .B(n22406), .C(n22405), .D(n22404), .Y(n34438)
         );
  AOI22XL U18169 ( .A0(n35130), .A1(n22403), .B0(n28465), .B1(n23089), .Y(
        n22404) );
  AOI22XL U18170 ( .A0(n34992), .A1(n22843), .B0(n26263), .B1(n22402), .Y(
        n22405) );
  AOI2BB1XL U18171 ( .A0N(n22401), .A1N(n35239), .B0(n22400), .Y(n22407) );
  INVXL U18172 ( .A(n23731), .Y(n35610) );
  AOI2BB1XL U18173 ( .A0N(conv_3[70]), .A1N(n31430), .B0(n31431), .Y(n32552)
         );
  AOI21XL U18174 ( .A0(n31478), .A1(n31473), .B0(n32163), .Y(n31430) );
  OAI2BB1XL U18175 ( .A0N(n32168), .A1N(n29676), .B0(n25246), .Y(n32606) );
  INVXL U18176 ( .A(n32606), .Y(n35598) );
  NOR2X1 U18177 ( .A(n32179), .B(n32177), .Y(n33823) );
  INVXL U18178 ( .A(n33818), .Y(n34392) );
  AOI22XL U18179 ( .A0(n34954), .A1(n22448), .B0(n23785), .B1(n22447), .Y(
        n22452) );
  OAI2BB1XL U18180 ( .A0N(n32184), .A1N(n29676), .B0(n25246), .Y(n33818) );
  AOI2BB1XL U18181 ( .A0N(conv_3[39]), .A1N(n31226), .B0(n35591), .Y(n31232)
         );
  AOI2BB1XL U18182 ( .A0N(conv_3[38]), .A1N(n35589), .B0(n35591), .Y(n31226)
         );
  OAI2BB1XL U18183 ( .A0N(n31303), .A1N(n29676), .B0(n25246), .Y(n33444) );
  INVXL U18184 ( .A(n33449), .Y(n35591) );
  AOI22XL U18185 ( .A0(N18471), .A1(n23786), .B0(n23785), .B1(n23784), .Y(
        n23787) );
  NOR2BXL U18186 ( .AN(n35577), .B(conv_3[26]), .Y(n35579) );
  AOI21XL U18187 ( .A0(conv_3[21]), .A1(n31274), .B0(n33002), .Y(n31262) );
  NOR2X1 U18188 ( .A(n33002), .B(n31274), .Y(n31273) );
  AOI21XL U18189 ( .A0(n31309), .A1(n29676), .B0(n18856), .Y(n35576) );
  AND2XL U18190 ( .A(n28640), .B(n28639), .Y(n32997) );
  INVXL U18191 ( .A(n27508), .Y(n34383) );
  NAND2X1 U18192 ( .A(n19229), .B(n19246), .Y(n19227) );
  NAND4XL U18193 ( .A(n18190), .B(n36247), .C(n18189), .D(n18188), .Y(n19185)
         );
  INVX2 U18194 ( .A(n18174), .Y(n19004) );
  AOI22XL U18195 ( .A0(n36246), .A1(n22525), .B0(n22522), .B1(n22713), .Y(
        n21661) );
  AOI22XL U18196 ( .A0(n36246), .A1(n22578), .B0(n22579), .B1(n22765), .Y(
        n21600) );
  AOI22XL U18197 ( .A0(n25299), .A1(conv_1[276]), .B0(n22615), .B1(conv_1[321]), .Y(n19944) );
  AOI22XL U18198 ( .A0(n25306), .A1(conv_1[112]), .B0(n22615), .B1(conv_1[142]), .Y(n19993) );
  AOI22XL U18199 ( .A0(n25306), .A1(conv_1[52]), .B0(n16662), .B1(conv_1[67]), 
        .Y(n19995) );
  AOI22XL U18200 ( .A0(n25306), .A1(conv_1[292]), .B0(n16673), .B1(conv_1[322]), .Y(n19998) );
  NOR2X1 U18201 ( .A(n22717), .B(n26796), .Y(n19899) );
  AOI22XL U18202 ( .A0(n36246), .A1(n22521), .B0(n22522), .B1(n22765), .Y(
        n21657) );
  AOI22XL U18203 ( .A0(n25306), .A1(conv_1[293]), .B0(n22690), .B1(conv_1[278]), .Y(n19978) );
  AOI22XL U18204 ( .A0(n16662), .A1(conv_1[308]), .B0(n22615), .B1(conv_1[323]), .Y(n19979) );
  AOI22XL U18205 ( .A0(n25306), .A1(conv_1[53]), .B0(n16662), .B1(conv_1[68]), 
        .Y(n19972) );
  AOI22XL U18206 ( .A0(n25299), .A1(conv_1[38]), .B0(n22615), .B1(conv_1[83]), 
        .Y(n19973) );
  AOI22XL U18207 ( .A0(n25306), .A1(conv_1[353]), .B0(n22615), .B1(conv_1[383]), .Y(n19974) );
  AOI22XL U18208 ( .A0(n36246), .A1(n22555), .B0(n22556), .B1(n22765), .Y(
        n21623) );
  AOI22XL U18209 ( .A0(n16662), .A1(conv_2[311]), .B0(n22615), .B1(conv_2[326]), .Y(n20894) );
  AOI22XL U18210 ( .A0(n16666), .A1(conv_2[356]), .B0(n22615), .B1(conv_2[386]), .Y(n20900) );
  AOI22XL U18211 ( .A0(n36246), .A1(n20946), .B0(n25915), .B1(n21358), .Y(
        n25917) );
  AOI22XL U18212 ( .A0(n22770), .A1(conv_2[351]), .B0(n22615), .B1(conv_2[381]), .Y(n20913) );
  AOI22XL U18213 ( .A0(n25299), .A1(conv_2[96]), .B0(n22615), .B1(conv_2[141]), 
        .Y(n20911) );
  AOI22XL U18214 ( .A0(n16662), .A1(conv_2[185]), .B0(n22615), .B1(conv_2[200]), .Y(n20822) );
  AOI22XL U18215 ( .A0(n16662), .A1(conv_2[305]), .B0(n22615), .B1(conv_2[320]), .Y(n20826) );
  AOI22XL U18216 ( .A0(n25299), .A1(conv_2[95]), .B0(n22615), .B1(conv_2[140]), 
        .Y(n20824) );
  AOI22XL U18217 ( .A0(n22770), .A1(conv_2[50]), .B0(n22615), .B1(conv_2[80]), 
        .Y(n20829) );
  AOI22XL U18218 ( .A0(n16662), .A1(conv_2[368]), .B0(n22615), .B1(conv_2[383]), .Y(n20795) );
  AOI22XL U18219 ( .A0(n22690), .A1(conv_2[278]), .B0(n22615), .B1(conv_2[323]), .Y(n20802) );
  NAND2XL U18220 ( .A(n36246), .B(n20878), .Y(n25989) );
  NAND2XL U18221 ( .A(n36246), .B(n21914), .Y(n26037) );
  AOI22XL U18222 ( .A0(n25289), .A1(conv_2[401]), .B0(n22690), .B1(conv_2[371]), .Y(n18330) );
  AOI22XL U18223 ( .A0(n16666), .A1(conv_3[175]), .B0(n25289), .B1(conv_3[190]), .Y(n19430) );
  AOI22XL U18224 ( .A0(n22759), .A1(conv_3[160]), .B0(n22615), .B1(conv_3[205]), .Y(n19431) );
  AOI22XL U18225 ( .A0(n16666), .A1(conv_3[55]), .B0(n22615), .B1(conv_3[85]), 
        .Y(n19442) );
  AOI211XL U18226 ( .A0(conv_3[200]), .A1(n22615), .B0(n19282), .C0(n19281), 
        .Y(n21244) );
  AOI22XL U18227 ( .A0(n25299), .A1(conv_3[276]), .B0(n22615), .B1(conv_3[321]), .Y(n19328) );
  AOI22XL U18228 ( .A0(n22759), .A1(conv_3[336]), .B0(n22615), .B1(conv_3[381]), .Y(n19322) );
  AOI211XL U18229 ( .A0(conv_3[308]), .A1(n25289), .B0(n19403), .C0(n19402), 
        .Y(n21339) );
  AOI22XL U18230 ( .A0(n16666), .A1(conv_3[295]), .B0(n25289), .B1(conv_3[310]), .Y(n19432) );
  AOI22XL U18231 ( .A0(n36246), .A1(n21359), .B0(n21357), .B1(n22765), .Y(
        n21363) );
  NOR2X1 U18232 ( .A(n22550), .B(n31435), .Y(n18513) );
  NOR2X1 U18233 ( .A(n18750), .B(n29166), .Y(n18518) );
  INVXL U18234 ( .A(n17749), .Y(n17850) );
  NOR4XL U18235 ( .A(n17118), .B(n17117), .C(n17116), .D(n17115), .Y(n17150)
         );
  NOR4XL U18236 ( .A(n17138), .B(n17137), .C(n17136), .D(n17135), .Y(n17149)
         );
  NOR2X1 U18237 ( .A(n21810), .B(n23053), .Y(n17799) );
  NOR2X1 U18238 ( .A(n22717), .B(n35239), .Y(n17896) );
  NOR2X1 U18239 ( .A(n19902), .B(n26274), .Y(n17790) );
  NAND2XL U18240 ( .A(n17923), .B(n18516), .Y(n17973) );
  INVXL U18241 ( .A(n17922), .Y(n18151) );
  INVXL U18242 ( .A(n17940), .Y(n18149) );
  INVXL U18243 ( .A(n17943), .Y(n18147) );
  INVXL U18244 ( .A(n18118), .Y(n18108) );
  INVXL U18245 ( .A(n17946), .Y(n18145) );
  NAND2XL U18246 ( .A(n36246), .B(n22471), .Y(n21564) );
  AOI22XL U18247 ( .A0(n25306), .A1(conv_1[172]), .B0(n16673), .B1(conv_1[202]), .Y(n19996) );
  NAND2XL U18248 ( .A(n36246), .B(n22623), .Y(n21581) );
  AOI22XL U18249 ( .A0(n25306), .A1(conv_1[173]), .B0(n22616), .B1(conv_1[158]), .Y(n19976) );
  AOI22XL U18250 ( .A0(n16662), .A1(conv_1[188]), .B0(n22615), .B1(conv_1[203]), .Y(n19977) );
  AOI211XL U18251 ( .A0(conv_1[130]), .A1(n25289), .B0(n19920), .C0(n19919), 
        .Y(n21636) );
  NAND2XL U18252 ( .A(n36246), .B(n22463), .Y(n21566) );
  AOI22XL U18253 ( .A0(n16662), .A1(conv_1[126]), .B0(n22615), .B1(conv_1[141]), .Y(n19939) );
  AOI22XL U18254 ( .A0(n22759), .A1(conv_1[156]), .B0(n22615), .B1(conv_1[201]), .Y(n19942) );
  OAI211XL U18255 ( .A0(n36246), .A1(n22560), .B0(n28528), .C0(n20274), .Y(
        n20275) );
  NAND2XL U18256 ( .A(n36246), .B(n22555), .Y(n20274) );
  AOI22XL U18257 ( .A0(n25306), .A1(conv_1[113]), .B0(n22615), .B1(conv_1[143]), .Y(n19970) );
  NOR2X1 U18258 ( .A(n22489), .B(n26026), .Y(n20293) );
  AOI22XL U18259 ( .A0(n25306), .A1(conv_1[118]), .B0(n16662), .B1(conv_1[133]), .Y(n20047) );
  AOI22XL U18260 ( .A0(n34963), .A1(n21610), .B0(n21600), .B1(n24056), .Y(
        n20026) );
  AOI22XL U18261 ( .A0(n28528), .A1(n21580), .B0(n34963), .B1(n21585), .Y(
        n20004) );
  AOI22XL U18262 ( .A0(n34963), .A1(n21627), .B0(n35234), .B1(n21624), .Y(
        n19982) );
  AOI2BB2XL U18263 ( .B0(n30029), .B1(n18526), .A0N(n19855), .A1N(conv_1[476]), 
        .Y(n22590) );
  NOR2X1 U18264 ( .A(n28488), .B(n26274), .Y(n25329) );
  AOI22XL U18265 ( .A0(n25306), .A1(conv_1[384]), .B0(n22690), .B1(conv_1[369]), .Y(n22531) );
  AOI22XL U18266 ( .A0(n25306), .A1(conv_1[324]), .B0(n16662), .B1(conv_1[339]), .Y(n22536) );
  AOI22XL U18267 ( .A0(n34963), .A1(n28473), .B0(n26585), .B1(n26451), .Y(
        n26428) );
  AOI22XL U18268 ( .A0(n36246), .A1(n22579), .B0(n22578), .B1(n21358), .Y(
        n28494) );
  AOI22XL U18269 ( .A0(n34963), .A1(n26595), .B0(n16663), .B1(n26594), .Y(
        n26596) );
  AOI22XL U18270 ( .A0(n36246), .A1(n22489), .B0(n22488), .B1(n22765), .Y(
        n28450) );
  AOI22XL U18271 ( .A0(n25306), .A1(conv_1[144]), .B0(n16662), .B1(conv_1[159]), .Y(n22533) );
  AOI22XL U18272 ( .A0(n25306), .A1(conv_1[203]), .B0(n16662), .B1(conv_1[218]), .Y(n22559) );
  AOI22XL U18273 ( .A0(n25306), .A1(conv_1[84]), .B0(n16662), .B1(conv_1[99]), 
        .Y(n22528) );
  AOI211XL U18274 ( .A0(conv_1[85]), .A1(n25306), .B0(n22492), .C0(n22491), 
        .Y(n28457) );
  AOI22XL U18275 ( .A0(n25306), .A1(conv_1[145]), .B0(n16673), .B1(conv_1[175]), .Y(n22480) );
  AOI211XL U18276 ( .A0(conv_1[96]), .A1(n25289), .B0(n22466), .C0(n22465), 
        .Y(n28505) );
  NOR2X1 U18277 ( .A(n22717), .B(n27105), .Y(n22466) );
  AOI22XL U18278 ( .A0(n36246), .A1(n22556), .B0(n22555), .B1(n21358), .Y(
        n28436) );
  NOR2X1 U18279 ( .A(n22457), .B(n22456), .Y(n28500) );
  NOR2X1 U18280 ( .A(n22612), .B(n35436), .Y(n22552) );
  AOI22XL U18281 ( .A0(n25306), .A1(conv_1[320]), .B0(n22616), .B1(conv_1[305]), .Y(n22566) );
  AOI22XL U18282 ( .A0(n25306), .A1(conv_1[380]), .B0(n16662), .B1(conv_1[395]), .Y(n22575) );
  AOI22XL U18283 ( .A0(n36246), .A1(n22522), .B0(n22521), .B1(n22743), .Y(
        n28517) );
  AOI22XL U18284 ( .A0(n25306), .A1(conv_1[24]), .B0(n16662), .B1(conv_1[39]), 
        .Y(n22526) );
  NOR2X1 U18285 ( .A(n22550), .B(n25287), .Y(n22482) );
  AOI211XL U18286 ( .A0(conv_1[235]), .A1(n22615), .B0(n22484), .C0(n22483), 
        .Y(n28456) );
  NOR2X1 U18287 ( .A(n22612), .B(n23295), .Y(n22484) );
  NOR2X1 U18288 ( .A(n22717), .B(n23155), .Y(n22478) );
  AOI211XL U18289 ( .A0(n22759), .A1(conv_1[10]), .B0(n22486), .C0(n22485), 
        .Y(n28463) );
  AOI211XL U18290 ( .A0(conv_2[370]), .A1(n25289), .B0(n20854), .C0(n20853), 
        .Y(n26040) );
  NAND2XL U18291 ( .A(n36246), .B(n26065), .Y(n21046) );
  AOI22XL U18292 ( .A0(n21011), .A1(conv_2[350]), .B0(n25289), .B1(conv_2[365]), .Y(n20820) );
  AOI22XL U18293 ( .A0(n25299), .A1(conv_2[335]), .B0(n22615), .B1(conv_2[380]), .Y(n20819) );
  AOI22XL U18294 ( .A0(n16662), .A1(conv_2[306]), .B0(n22615), .B1(conv_2[321]), .Y(n20918) );
  AOI22XL U18295 ( .A0(n16662), .A1(conv_2[188]), .B0(n22615), .B1(conv_2[203]), .Y(n20797) );
  NOR2X1 U18296 ( .A(n25977), .B(n20810), .Y(n25974) );
  AOI22XL U18297 ( .A0(n36246), .A1(n25988), .B0(n25997), .B1(n21358), .Y(
        n25993) );
  AOI22XL U18298 ( .A0(n25306), .A1(conv_2[57]), .B0(n16662), .B1(conv_2[72]), 
        .Y(n21043) );
  AOI22XL U18299 ( .A0(n22690), .A1(conv_2[42]), .B0(n22615), .B1(conv_2[87]), 
        .Y(n21042) );
  AOI22XL U18300 ( .A0(n25306), .A1(conv_2[177]), .B0(n25289), .B1(conv_2[192]), .Y(n21045) );
  AOI22XL U18301 ( .A0(n22690), .A1(conv_2[162]), .B0(n22615), .B1(conv_2[207]), .Y(n21044) );
  AOI22XL U18302 ( .A0(n34963), .A1(n25920), .B0(n24056), .B1(n25917), .Y(
        n21907) );
  AOI22XL U18303 ( .A0(n36246), .A1(n25958), .B0(n25955), .B1(n22743), .Y(
        n25956) );
  AOI2BB2XL U18304 ( .B0(n34963), .B1(n25903), .A0N(n19767), .A1N(n25896), .Y(
        n21881) );
  AOI22XL U18305 ( .A0(n16659), .A1(n25984), .B0(n34963), .B1(n25978), .Y(
        n21934) );
  AOI22XL U18306 ( .A0(n34963), .A1(n26018), .B0(n26015), .B1(n24056), .Y(
        n21928) );
  AOI22XL U18307 ( .A0(n22690), .A1(conv_2[280]), .B0(n22615), .B1(conv_2[325]), .Y(n20849) );
  AOI22XL U18308 ( .A0(n22770), .A1(conv_2[175]), .B0(n22615), .B1(conv_2[205]), .Y(n20846) );
  NOR2X1 U18309 ( .A(n18271), .B(n18270), .Y(n25176) );
  AOI22XL U18310 ( .A0(n36246), .A1(n21913), .B0(n21914), .B1(n21688), .Y(
        n25586) );
  AOI22XL U18311 ( .A0(n25289), .A1(conv_2[337]), .B0(n16673), .B1(conv_2[352]), .Y(n18300) );
  AOI22XL U18312 ( .A0(n25289), .A1(conv_2[335]), .B0(n22690), .B1(conv_2[305]), .Y(n18233) );
  AOI22XL U18313 ( .A0(n25289), .A1(conv_2[40]), .B0(n18658), .B1(conv_2[10]), 
        .Y(n18223) );
  AOI22XL U18314 ( .A0(n25289), .A1(conv_2[338]), .B0(n16673), .B1(conv_2[353]), .Y(n18315) );
  AOI22XL U18315 ( .A0(n25289), .A1(conv_2[398]), .B0(n22759), .B1(conv_2[368]), .Y(n18313) );
  AOI22XL U18316 ( .A0(n36246), .A1(n20803), .B0(n21931), .B1(n22743), .Y(
        n25560) );
  AOI22XL U18317 ( .A0(n36246), .A1(n26027), .B0(n26009), .B1(n22743), .Y(
        n25156) );
  AOI22XL U18318 ( .A0(n36246), .A1(n25997), .B0(n25988), .B1(n21688), .Y(
        n25174) );
  AOI211XL U18319 ( .A0(n25289), .A1(conv_2[215]), .B0(n18230), .C0(n18229), 
        .Y(n25141) );
  AOI22XL U18320 ( .A0(n25289), .A1(conv_2[159]), .B0(n16673), .B1(conv_2[174]), .Y(n18268) );
  AOI2BB2XL U18321 ( .B0(n36245), .B1(n25570), .A0N(n25576), .A1N(n36245), .Y(
        n24766) );
  AOI22XL U18322 ( .A0(n25289), .A1(conv_2[158]), .B0(n16673), .B1(conv_2[173]), .Y(n18318) );
  AOI211XL U18323 ( .A0(n25289), .A1(conv_2[216]), .B0(n18292), .C0(n18291), 
        .Y(n25543) );
  AOI22XL U18324 ( .A0(n25289), .A1(conv_2[341]), .B0(n22690), .B1(conv_2[311]), .Y(n18333) );
  AOI22XL U18325 ( .A0(n25289), .A1(conv_2[340]), .B0(n22759), .B1(conv_2[310]), .Y(n18216) );
  AOI22XL U18326 ( .A0(n25289), .A1(conv_2[400]), .B0(n22690), .B1(conv_2[370]), .Y(n18214) );
  AOI211XL U18327 ( .A0(conv_2[160]), .A1(n25289), .B0(n18220), .C0(n18219), 
        .Y(n25597) );
  AOI211XL U18328 ( .A0(conv_2[218]), .A1(n25289), .B0(n18323), .C0(n18322), 
        .Y(n25566) );
  AOI22XL U18329 ( .A0(n25289), .A1(conv_2[38]), .B0(n22690), .B1(conv_2[8]), 
        .Y(n18319) );
  NOR2X1 U18330 ( .A(n20563), .B(n22713), .Y(n21425) );
  AOI22XL U18331 ( .A0(n16666), .A1(conv_3[352]), .B0(n22615), .B1(conv_3[382]), .Y(n19394) );
  AOI22XL U18332 ( .A0(n16662), .A1(conv_3[67]), .B0(n22615), .B1(conv_3[82]), 
        .Y(n19385) );
  NOR2X1 U18333 ( .A(n22612), .B(n33835), .Y(n19429) );
  AOI211XL U18334 ( .A0(conv_3[115]), .A1(n25306), .B0(n19426), .C0(n19425), 
        .Y(n21356) );
  AOI22XL U18335 ( .A0(n22759), .A1(conv_3[279]), .B0(n22615), .B1(conv_3[324]), .Y(n19338) );
  AOI22XL U18336 ( .A0(n16666), .A1(conv_3[174]), .B0(n25289), .B1(conv_3[189]), .Y(n19336) );
  AOI22XL U18337 ( .A0(n22759), .A1(conv_3[159]), .B0(n22615), .B1(conv_3[204]), .Y(n19337) );
  AOI22XL U18338 ( .A0(n36246), .A1(n21286), .B0(n21295), .B1(n22743), .Y(
        n21289) );
  NOR2X1 U18339 ( .A(n22550), .B(n31969), .Y(n19302) );
  NOR2X1 U18340 ( .A(n19579), .B(n19578), .Y(n21407) );
  AOI22XL U18341 ( .A0(n16666), .A1(conv_3[298]), .B0(n22615), .B1(conv_3[328]), .Y(n19583) );
  NOR2X1 U18342 ( .A(n20562), .B(n21425), .Y(n21435) );
  AOI211XL U18343 ( .A0(conv_3[132]), .A1(n25289), .B0(n19546), .C0(n19545), 
        .Y(n21428) );
  AOI22XL U18344 ( .A0(n34963), .A1(n21229), .B0(n34961), .B1(n21212), .Y(
        n20466) );
  AOI22XL U18345 ( .A0(n36246), .A1(n21213), .B0(n21226), .B1(n22713), .Y(
        n21216) );
  AOI22XL U18346 ( .A0(n16662), .A1(conv_3[126]), .B0(n22615), .B1(conv_3[141]), .Y(n19320) );
  AOI22XL U18347 ( .A0(n16667), .A1(n21266), .B0(n34963), .B1(n21271), .Y(
        n20456) );
  AOI22XL U18348 ( .A0(n36246), .A1(n21269), .B0(n21263), .B1(n21688), .Y(
        n21262) );
  AOI22XL U18349 ( .A0(n34963), .A1(n21307), .B0(n34961), .B1(n21306), .Y(
        n20480) );
  AOI22XL U18350 ( .A0(n25306), .A1(conv_3[324]), .B0(n22615), .B1(conv_3[354]), .Y(n18567) );
  AOI22XL U18351 ( .A0(n22762), .A1(conv_3[321]), .B0(n22615), .B1(conv_3[351]), .Y(n18550) );
  AOI22XL U18352 ( .A0(n18658), .A1(conv_3[366]), .B0(n22615), .B1(conv_3[411]), .Y(n18544) );
  AOI22XL U18353 ( .A0(n16659), .A1(n26232), .B0(n34963), .B1(n35116), .Y(
        n18590) );
  NOR2X1 U18354 ( .A(n16668), .B(n31619), .Y(n18460) );
  AOI22XL U18355 ( .A0(n25306), .A1(conv_3[144]), .B0(n16662), .B1(conv_3[159]), .Y(n18570) );
  NOR2X1 U18356 ( .A(n22550), .B(n31595), .Y(n18474) );
  AOI211XL U18357 ( .A0(n22616), .A1(conv_3[10]), .B0(n18515), .C0(n18514), 
        .Y(n35055) );
  AOI22XL U18358 ( .A0(n16662), .A1(conv_3[96]), .B0(n22615), .B1(conv_3[111]), 
        .Y(n18548) );
  AOI22XL U18359 ( .A0(n18658), .A1(conv_3[365]), .B0(n22615), .B1(conv_3[410]), .Y(n18457) );
  AOI22XL U18360 ( .A0(n16666), .A1(conv_3[20]), .B0(n22615), .B1(conv_3[50]), 
        .Y(n18454) );
  AOI22XL U18361 ( .A0(n16666), .A1(conv_3[80]), .B0(n22615), .B1(conv_3[110]), 
        .Y(n18465) );
  AOI22XL U18362 ( .A0(n36246), .A1(n21242), .B0(n21236), .B1(n22713), .Y(
        n35045) );
  AOI22XL U18363 ( .A0(n36246), .A1(n20513), .B0(n20514), .B1(n22743), .Y(
        n35034) );
  AOI22XL U18364 ( .A0(n16666), .A1(conv_3[325]), .B0(n25289), .B1(conv_3[340]), .Y(n18508) );
  AOI22XL U18365 ( .A0(n36246), .A1(n21357), .B0(n21359), .B1(n21688), .Y(
        n35054) );
  AOI22XL U18366 ( .A0(n36246), .A1(n21295), .B0(n21286), .B1(n22743), .Y(
        n35081) );
  INVXL U18367 ( .A(n22368), .Y(n18777) );
  NOR2X1 U18368 ( .A(n21944), .B(n17172), .Y(n17853) );
  NOR2X1 U18369 ( .A(n17171), .B(n19182), .Y(n17843) );
  NOR2X1 U18370 ( .A(n28467), .B(n19182), .Y(n17841) );
  NOR2X1 U18371 ( .A(n16669), .B(n17172), .Y(n17754) );
  INVXL U18372 ( .A(n17848), .Y(n17690) );
  NOR2X1 U18373 ( .A(n16760), .B(n21944), .Y(n17787) );
  NOR2X1 U18374 ( .A(n19902), .B(n26621), .Y(n17816) );
  NOR2X1 U18375 ( .A(n20755), .B(n18119), .Y(n17822) );
  NOR2X1 U18376 ( .A(n34969), .B(n20726), .Y(n17900) );
  NAND4XL U18377 ( .A(n17436), .B(n17435), .C(n17434), .D(n17433), .Y(n17437)
         );
  INVXL U18378 ( .A(n17166), .Y(n17172) );
  INVXL U18379 ( .A(n17748), .Y(n17851) );
  NOR2X1 U18380 ( .A(n17170), .B(n17172), .Y(n17752) );
  ADDFXL U18381 ( .A(n17509), .B(affine_1[17]), .CI(n17508), .CO(
        DP_OP_5167J1_123_9881_n18), .S(DP_OP_5167J1_123_9881_n19) );
  AND2XL U18382 ( .A(n17161), .B(n17918), .Y(DP_OP_5166J1_122_9881_n60) );
  NAND2XL U18383 ( .A(n16734), .B(n17169), .Y(n17746) );
  INVXL U18384 ( .A(n17747), .Y(n17852) );
  INVXL U18385 ( .A(n17753), .Y(n17837) );
  NOR2X1 U18386 ( .A(n16760), .B(n16669), .Y(n17798) );
  NOR2X1 U18387 ( .A(n21944), .B(n23053), .Y(n17883) );
  NOR2X1 U18388 ( .A(n19416), .B(n23053), .Y(n17865) );
  NOR2X1 U18389 ( .A(n26207), .B(n18118), .Y(n17804) );
  NOR2X1 U18390 ( .A(n20755), .B(n18116), .Y(n17887) );
  NOR2X1 U18391 ( .A(n26207), .B(n18117), .Y(n17898) );
  AND2XL U18392 ( .A(n19097), .B(n23785), .Y(n17803) );
  NOR2X1 U18393 ( .A(n22550), .B(n26279), .Y(n17868) );
  NOR2X1 U18394 ( .A(n17170), .B(n23052), .Y(n17800) );
  NOR2X1 U18395 ( .A(n20726), .B(n25853), .Y(n17875) );
  NOR2X1 U18396 ( .A(n17170), .B(n26409), .Y(n17797) );
  NOR2X1 U18397 ( .A(n16669), .B(n23053), .Y(n17791) );
  NOR2X1 U18398 ( .A(n26207), .B(n18109), .Y(n17878) );
  NOR2X1 U18399 ( .A(n34969), .B(n17165), .Y(n17877) );
  NOR2X1 U18400 ( .A(n34989), .B(n21953), .Y(n17823) );
  NOR2X1 U18401 ( .A(n22550), .B(n26274), .Y(n16724) );
  NOR2X1 U18402 ( .A(n34969), .B(n17173), .Y(n17802) );
  NOR2X1 U18403 ( .A(n18750), .B(n28479), .Y(n17789) );
  NOR2X1 U18404 ( .A(n26207), .B(n18116), .Y(n17884) );
  NOR2X1 U18405 ( .A(n20755), .B(n18118), .Y(n17792) );
  NOR2X1 U18406 ( .A(n17170), .B(n23053), .Y(n17885) );
  NOR2X1 U18407 ( .A(n26207), .B(n18120), .Y(n17824) );
  NOR2X1 U18408 ( .A(n35135), .B(n22018), .Y(n17821) );
  NOR2X1 U18409 ( .A(n26207), .B(n18127), .Y(n17811) );
  NOR2X1 U18410 ( .A(n20755), .B(n18117), .Y(n17876) );
  ADDFXL U18411 ( .A(n17164), .B(affine_1[27]), .CI(n17163), .CO(
        DP_OP_5166J1_122_9881_n18), .S(DP_OP_5166J1_122_9881_n19) );
  INVXL U18412 ( .A(n18116), .Y(n18072) );
  AOI21XL U18413 ( .A0(n19221), .A1(n21830), .B0(n17923), .Y(n17972) );
  OAI211XL U18414 ( .A0(n20397), .A1(n18127), .B0(n18100), .C0(n18099), .Y(
        n19695) );
  NOR3XL U18415 ( .A(n18098), .B(n18097), .C(n18096), .Y(n18099) );
  OAI2BB1XL U18416 ( .A0N(weight_2[50]), .A1N(n18049), .B0(n18031), .Y(n19611)
         );
  MXI2XL U18417 ( .A(n24560), .B(n24561), .S0(n19694), .Y(n18059) );
  MXI2XL U18418 ( .A(n24560), .B(n24561), .S0(n19666), .Y(n18057) );
  AOI2BB2XL U18419 ( .B0(n20735), .B1(n30792), .A0N(conv_3[451]), .A1N(n35269), 
        .Y(n21144) );
  AOI2BB2XL U18420 ( .B0(n20735), .B1(n30597), .A0N(conv_3[241]), .A1N(n35269), 
        .Y(n21150) );
  OR2XL U18421 ( .A(n19147), .B(n23820), .Y(n19148) );
  NOR2X1 U18422 ( .A(n35272), .B(n23816), .Y(n19147) );
  NOR2X1 U18423 ( .A(n19127), .B(n23941), .Y(n19128) );
  NOR2X1 U18424 ( .A(n19125), .B(n33501), .Y(n19127) );
  NOR2X1 U18425 ( .A(n25072), .B(n33433), .Y(n25074) );
  NAND2XL U18426 ( .A(n36246), .B(n25854), .Y(n20983) );
  NOR2X1 U18427 ( .A(n36244), .B(n25119), .Y(n25125) );
  NOR2X1 U18428 ( .A(n23790), .B(n33987), .Y(n23792) );
  NOR2X1 U18429 ( .A(n19471), .B(n21830), .Y(n19474) );
  OAI21XL U18430 ( .A0(conv_3[496]), .A1(n30729), .B0(n30730), .Y(n27621) );
  NOR2X1 U18431 ( .A(n23202), .B(n23742), .Y(n23203) );
  NOR2X1 U18432 ( .A(n23199), .B(n23201), .Y(n23202) );
  AOI2BB2XL U18433 ( .B0(n20735), .B1(n23472), .A0N(conv_1[243]), .A1N(n35269), 
        .Y(n22638) );
  AND2XL U18434 ( .A(n22417), .B(n27020), .Y(n22418) );
  AOI222XL U18435 ( .A0(n27445), .A1(conv_1[17]), .B0(n27445), .B1(n27444), 
        .C0(conv_1[17]), .C1(n27444), .Y(n26501) );
  NAND2XL U18436 ( .A(n36246), .B(n25836), .Y(n25831) );
  AOI2BB1XL U18437 ( .A0N(n30323), .A1N(n30318), .B0(n30319), .Y(n18932) );
  AOI22XL U18438 ( .A0(n36246), .A1(n21123), .B0(n20422), .B1(n21358), .Y(
        n21132) );
  NOR2X1 U18439 ( .A(n25698), .B(n28292), .Y(n35129) );
  AOI2BB2XL U18440 ( .B0(n20735), .B1(n30189), .A0N(conv_3[453]), .A1N(n35269), 
        .Y(n21124) );
  OAI21XL U18441 ( .A0(conv_3[497]), .A1(n30723), .B0(n30724), .Y(n27623) );
  AOI222XL U18442 ( .A0(n30818), .A1(conv_3[152]), .B0(n30818), .B1(n30817), 
        .C0(conv_3[152]), .C1(n30817), .Y(n22180) );
  NOR2XL U18443 ( .A(n29426), .B(n31418), .Y(n23898) );
  AOI22XL U18444 ( .A0(n25289), .A1(conv_1[184]), .B0(n22690), .B1(conv_1[154]), .Y(n19884) );
  AOI22XL U18445 ( .A0(n25289), .A1(conv_1[124]), .B0(n22690), .B1(conv_1[94]), 
        .Y(n19881) );
  AOI22XL U18446 ( .A0(n25289), .A1(conv_1[304]), .B0(n16673), .B1(conv_1[319]), .Y(n19883) );
  AOI2BB1XL U18447 ( .A0N(conv_1[438]), .A1N(n26939), .B0(n26940), .Y(n23641)
         );
  NOR2X1 U18448 ( .A(n35498), .B(n28070), .Y(n25252) );
  AOI222XL U18449 ( .A0(n23194), .A1(n23193), .B0(n23194), .B1(conv_1[378]), 
        .C0(n23193), .C1(conv_1[378]), .Y(n19150) );
  NOR2X1 U18450 ( .A(n35500), .B(n27532), .Y(n19152) );
  AOI2BB1XL U18451 ( .A0N(conv_1[198]), .A1N(n23539), .B0(n23540), .Y(n23437)
         );
  AOI2BB1XL U18452 ( .A0N(conv_1[183]), .A1N(n23611), .B0(n23612), .Y(n23590)
         );
  NOR2X1 U18453 ( .A(n35500), .B(n34703), .Y(n23591) );
  NOR2X1 U18454 ( .A(n35500), .B(n28948), .Y(n23649) );
  NOR2X1 U18455 ( .A(n35500), .B(n26509), .Y(n26513) );
  NOR2X1 U18456 ( .A(n35500), .B(n33988), .Y(n25078) );
  NOR2X1 U18457 ( .A(n21858), .B(n22014), .Y(n21860) );
  INVX4 U18458 ( .A(N17631), .Y(n18516) );
  AOI22XL U18459 ( .A0(n22762), .A1(conv_2[169]), .B0(n22615), .B1(conv_2[199]), .Y(n20786) );
  AOI222XL U18460 ( .A0(n29644), .A1(n29645), .B0(n29644), .B1(conv_2[513]), 
        .C0(n29645), .C1(conv_2[513]), .Y(n27767) );
  OAI2BB1XL U18461 ( .A0N(n34104), .A1N(n34099), .B0(n34100), .Y(n18933) );
  AOI2BB1XL U18462 ( .A0N(conv_2[483]), .A1N(n29547), .B0(n29548), .Y(n27739)
         );
  NOR2X1 U18463 ( .A(n27735), .B(n35858), .Y(n27740) );
  OAI21XL U18464 ( .A0(conv_2[468]), .A1(n29559), .B0(n29560), .Y(n27865) );
  AOI2BB1XL U18465 ( .A0N(conv_2[378]), .A1N(n23991), .B0(n23992), .Y(n23077)
         );
  AOI222XL U18466 ( .A0(n24185), .A1(conv_2[303]), .B0(n24185), .B1(n24184), 
        .C0(conv_2[303]), .C1(n24184), .Y(n19111) );
  NOR2X1 U18467 ( .A(n19108), .B(n35858), .Y(n19113) );
  NOR2X1 U18468 ( .A(n35858), .B(n31871), .Y(n28090) );
  NOR2X1 U18469 ( .A(n35858), .B(n34426), .Y(n22901) );
  NOR2X1 U18470 ( .A(n35858), .B(n28948), .Y(n23336) );
  AOI22XL U18471 ( .A0(n36246), .A1(n20492), .B0(n20495), .B1(n22765), .Y(
        n21191) );
  NOR2X1 U18472 ( .A(n20490), .B(n21960), .Y(n20494) );
  AOI22XL U18473 ( .A0(n36246), .A1(n20490), .B0(n20495), .B1(n21688), .Y(
        n21202) );
  AOI2BB1XL U18474 ( .A0N(conv_3[498]), .A1N(n29631), .B0(n29632), .Y(n27625)
         );
  NOR2X1 U18475 ( .A(n31691), .B(n33422), .Y(n27626) );
  AOI2BB1XL U18476 ( .A0N(conv_3[423]), .A1N(n31693), .B0(n31692), .Y(n31694)
         );
  AOI2BB1XL U18477 ( .A0N(conv_3[393]), .A1N(n29695), .B0(n29696), .Y(n23632)
         );
  NOR2X1 U18478 ( .A(n31691), .B(n32016), .Y(n23633) );
  NOR2X1 U18479 ( .A(n31691), .B(n23504), .Y(n23509) );
  OR2XL U18480 ( .A(n35565), .B(n35562), .Y(n23805) );
  NOR2X1 U18481 ( .A(n34703), .B(n31691), .Y(n22133) );
  OAI21XL U18482 ( .A0(conv_3[153]), .A1(n29959), .B0(n29960), .Y(n22182) );
  NOR2X1 U18483 ( .A(n31691), .B(n33020), .Y(n22921) );
  NAND2XL U18484 ( .A(n36246), .B(n22766), .Y(n21726) );
  AOI22XL U18485 ( .A0(n25306), .A1(conv_1[58]), .B0(n16662), .B1(conv_1[73]), 
        .Y(n20050) );
  NOR2X1 U18486 ( .A(n21616), .B(n21615), .Y(n21697) );
  NAND2XL U18487 ( .A(n36246), .B(n22720), .Y(n20194) );
  AOI22XL U18488 ( .A0(n28528), .A1(n21757), .B0(n34963), .B1(n21754), .Y(
        n20081) );
  AOI22XL U18489 ( .A0(n28528), .A1(n21734), .B0(n34963), .B1(n21727), .Y(
        n20054) );
  AOI22XL U18490 ( .A0(n36246), .A1(n22720), .B0(n22721), .B1(n22743), .Y(
        n21708) );
  AOI211XL U18491 ( .A0(conv_1[179]), .A1(n25306), .B0(n19771), .C0(n19770), 
        .Y(n21713) );
  NOR2X1 U18492 ( .A(n22740), .B(n32995), .Y(n19771) );
  AOI2BB2XL U18493 ( .B0(n34963), .B1(n21644), .A0N(n21637), .A1N(n35196), .Y(
        n19928) );
  AOI211XL U18494 ( .A0(n16667), .A1(n21679), .B0(n19968), .C0(n19967), .Y(
        n20040) );
  NOR2X1 U18495 ( .A(n33201), .B(n21953), .Y(n19859) );
  AOI22XL U18496 ( .A0(n34963), .A1(n28476), .B0(n26262), .B1(n28474), .Y(
        n25327) );
  NOR2X1 U18497 ( .A(n22707), .B(n22706), .Y(n28418) );
  AOI22XL U18498 ( .A0(n36246), .A1(n22767), .B0(n22766), .B1(n22765), .Y(
        n28550) );
  AOI211XL U18499 ( .A0(n26470), .A1(n26593), .B0(n26427), .C0(n26426), .Y(
        n26437) );
  AOI22XL U18500 ( .A0(n34963), .A1(n26586), .B0(n34984), .B1(n26588), .Y(
        n26424) );
  AOI22XL U18501 ( .A0(n16659), .A1(n28487), .B0(n34963), .B1(n28486), .Y(
        n26417) );
  AOI211XL U18502 ( .A0(n34963), .A1(n28529), .B0(n26446), .C0(n26445), .Y(
        n26447) );
  AOI22XL U18503 ( .A0(n34963), .A1(n26587), .B0(n28324), .B1(n26586), .Y(
        n26590) );
  AOI22XL U18504 ( .A0(n36246), .A1(n22745), .B0(n22744), .B1(n22743), .Y(
        n28570) );
  AOI211XL U18505 ( .A0(n25289), .A1(conv_1[43]), .B0(n22769), .C0(n22768), 
        .Y(n28552) );
  AOI222XL U18506 ( .A0(n35484), .A1(n35483), .B0(n35484), .B1(conv_1[409]), 
        .C0(n35483), .C1(conv_1[409]), .Y(n25253) );
  AOI222XL U18507 ( .A0(n30766), .A1(n30767), .B0(n30766), .B1(conv_1[274]), 
        .C0(n30767), .C1(conv_1[274]), .Y(n22287) );
  AOI22XL U18508 ( .A0(n19005), .A1(filter_1[12]), .B0(n16676), .B1(
        filter_1[36]), .Y(n18836) );
  AOI22XL U18509 ( .A0(filter_1[17]), .A1(n19005), .B0(filter_1[41]), .B1(
        n16676), .Y(n18726) );
  NOR2X1 U18510 ( .A(n35858), .B(n33429), .Y(n27687) );
  AOI22XL U18511 ( .A0(n25306), .A1(conv_2[357]), .B0(n16662), .B1(conv_2[372]), .Y(n21040) );
  AOI22XL U18512 ( .A0(n22759), .A1(conv_2[342]), .B0(n22615), .B1(conv_2[387]), .Y(n21039) );
  AOI211XL U18513 ( .A0(conv_2[133]), .A1(n25289), .B0(n21067), .C0(n21066), 
        .Y(n26088) );
  NOR2X1 U18514 ( .A(n26051), .B(n26054), .Y(n26050) );
  AOI22XL U18515 ( .A0(n28556), .A1(n26071), .B0(n34963), .B1(n26069), .Y(
        n22001) );
  AOI22XL U18516 ( .A0(n34963), .A1(n26093), .B0(n24056), .B1(n22022), .Y(
        n22023) );
  AOI211XL U18517 ( .A0(conv_2[134]), .A1(n25289), .B0(n20757), .C0(n20756), 
        .Y(n25821) );
  AOI211XL U18518 ( .A0(conv_2[179]), .A1(n25306), .B0(n20763), .C0(n20762), 
        .Y(n25823) );
  AOI211XL U18519 ( .A0(conv_2[374]), .A1(n25289), .B0(n20759), .C0(n20758), 
        .Y(n25820) );
  NOR2X1 U18520 ( .A(n16668), .B(n29453), .Y(n20759) );
  AOI22XL U18521 ( .A0(n34963), .A1(n25996), .B0(n34961), .B1(n25995), .Y(
        n21967) );
  NOR2X1 U18522 ( .A(n26002), .B(n22034), .Y(n22037) );
  NOR2X1 U18523 ( .A(n27919), .B(n21953), .Y(n21946) );
  AOI22XL U18524 ( .A0(n36246), .A1(n21997), .B0(n26065), .B1(n21358), .Y(
        n25636) );
  NOR2X1 U18525 ( .A(n25052), .B(n25048), .Y(n25026) );
  AOI22XL U18526 ( .A0(n34963), .A1(n25526), .B0(n16670), .B1(n25531), .Y(
        n24082) );
  AOI211XL U18527 ( .A0(n34963), .A1(n25601), .B0(n24067), .C0(n24066), .Y(
        n24068) );
  AOI22XL U18528 ( .A0(n34963), .A1(n25517), .B0(n25519), .B1(n28372), .Y(
        n24732) );
  AOI22XL U18529 ( .A0(n34963), .A1(n25530), .B0(n25147), .B1(n28372), .Y(
        n24736) );
  AOI211XL U18530 ( .A0(n34963), .A1(n24746), .B0(n24745), .C0(n24744), .Y(
        n24754) );
  AOI2BB2XL U18531 ( .B0(n36245), .B1(n25649), .A0N(n25653), .A1N(n36245), .Y(
        n24793) );
  NOR2X1 U18532 ( .A(n22612), .B(n33267), .Y(n18407) );
  AOI22XL U18533 ( .A0(n36246), .A1(n21059), .B0(n22012), .B1(n22743), .Y(
        n25652) );
  AOI22XL U18534 ( .A0(n25289), .A1(conv_2[44]), .B0(n16723), .B1(conv_2[59]), 
        .Y(n18200) );
  AOI22XL U18535 ( .A0(n25306), .A1(conv_2[88]), .B0(n25289), .B1(conv_2[103]), 
        .Y(n18416) );
  AOI22XL U18536 ( .A0(n36246), .A1(n25812), .B0(n21976), .B1(n22765), .Y(
        n25624) );
  AOI22XL U18537 ( .A0(n25289), .A1(conv_2[404]), .B0(n16723), .B1(conv_2[419]), .Y(n18193) );
  AOI2BB1XL U18538 ( .A0N(conv_2[499]), .A1N(n28989), .B0(n28990), .Y(n18935)
         );
  OAI21XL U18539 ( .A0(conv_2[469]), .A1(n28995), .B0(n28996), .Y(n27867) );
  AOI22XL U18540 ( .A0(n19007), .A1(filter_2[28]), .B0(n19005), .B1(
        filter_2[16]), .Y(n18905) );
  OAI21XL U18541 ( .A0(conv_2[364]), .A1(n23356), .B0(n23357), .Y(n23125) );
  OAI2BB1XL U18542 ( .A0N(n34407), .A1N(n34402), .B0(n34403), .Y(n25679) );
  NAND2XL U18543 ( .A(n30220), .B(n30939), .Y(n30204) );
  OAI2BB1XL U18544 ( .A0N(n25280), .A1N(n25275), .B0(n25276), .Y(n18971) );
  AOI22XL U18545 ( .A0(n19005), .A1(filter_2[12]), .B0(n16676), .B1(
        filter_2[36]), .Y(n18917) );
  AOI32XL U18546 ( .A0(n22343), .A1(n22342), .A2(n22341), .B0(n22716), .B1(
        n22342), .Y(n22344) );
  AOI211XL U18547 ( .A0(n22368), .A1(n22340), .B0(n22339), .C0(n22338), .Y(
        n22342) );
  AOI22XL U18548 ( .A0(n19005), .A1(filter_2[17]), .B0(n16676), .B1(
        filter_2[41]), .Y(n18898) );
  NOR2X1 U18549 ( .A(n31691), .B(n33429), .Y(n23550) );
  OR2XL U18550 ( .A(n36246), .B(n18196), .Y(n21237) );
  AOI211XL U18551 ( .A0(conv_3[192]), .A1(n25289), .B0(n19560), .C0(n19559), 
        .Y(n21430) );
  OR4XL U18552 ( .A(n21279), .B(n21278), .C(n21277), .D(n21276), .Y(n21374) );
  AOI31XL U18553 ( .A0(n36246), .A1(n16664), .A2(n21333), .B0(n21332), .Y(
        n21350) );
  NAND2XL U18554 ( .A(n36246), .B(n21403), .Y(n19575) );
  AOI211XL U18555 ( .A0(conv_3[73]), .A1(n25289), .B0(n19574), .C0(n19573), 
        .Y(n21408) );
  AOI22XL U18556 ( .A0(n16716), .A1(conv_3[193]), .B0(n22615), .B1(conv_3[208]), .Y(n19568) );
  NOR2X1 U18557 ( .A(n19424), .B(n19423), .Y(n19590) );
  AOI22XL U18558 ( .A0(n36246), .A1(n20554), .B0(n20553), .B1(n22765), .Y(
        n21409) );
  AOI22XL U18559 ( .A0(n22759), .A1(conv_3[103]), .B0(n22615), .B1(conv_3[148]), .Y(n19580) );
  NOR2X1 U18560 ( .A(n21944), .B(n32190), .Y(n19570) );
  NOR2X1 U18561 ( .A(n19524), .B(n19523), .Y(n21393) );
  NOR2X1 U18562 ( .A(n20542), .B(n21382), .Y(n21385) );
  AOI211XL U18563 ( .A0(conv_3[134]), .A1(n25289), .B0(n19528), .C0(n19527), 
        .Y(n21389) );
  AOI211XL U18564 ( .A0(conv_3[194]), .A1(n25289), .B0(n19526), .C0(n19525), 
        .Y(n21390) );
  AOI22XL U18565 ( .A0(n16666), .A1(conv_3[299]), .B0(n25289), .B1(conv_3[314]), .Y(n19534) );
  AOI22XL U18566 ( .A0(n22759), .A1(conv_3[284]), .B0(n22615), .B1(conv_3[329]), .Y(n19533) );
  AOI211XL U18567 ( .A0(n34963), .A1(n21241), .B0(n20505), .C0(n20504), .Y(
        n20510) );
  AOI22XL U18568 ( .A0(n34963), .A1(n21346), .B0(n35234), .B1(n21334), .Y(
        n20521) );
  OR2XL U18569 ( .A(n36246), .B(n26274), .Y(n22009) );
  INVXL U18570 ( .A(n19098), .Y(n17170) );
  INVXL U18571 ( .A(n19416), .Y(n21990) );
  INVX2 U18572 ( .A(n22014), .Y(n21991) );
  AOI211XL U18573 ( .A0(n34963), .A1(n35094), .B0(n26221), .C0(n26220), .Y(
        n26236) );
  AOI22XL U18574 ( .A0(n28528), .A1(n35115), .B0(n34963), .B1(n35123), .Y(
        n26234) );
  AOI22XL U18575 ( .A0(n16666), .A1(conv_3[387]), .B0(n22615), .B1(conv_3[417]), .Y(n18695) );
  AOI22XL U18576 ( .A0(n16667), .A1(n35185), .B0(n34963), .B1(n35179), .Y(
        n24877) );
  INVXL U18577 ( .A(n16673), .Y(n18321) );
  INVX2 U18578 ( .A(n18810), .Y(n22740) );
  AOI22XL U18579 ( .A0(n22347), .A1(conv_3[147]), .B0(n22615), .B1(conv_3[177]), .Y(n18693) );
  AOI22XL U18580 ( .A0(n36246), .A1(n19558), .B0(n20563), .B1(n21358), .Y(
        n35206) );
  INVX3 U18581 ( .A(n18321), .Y(n22615) );
  AOI22XL U18582 ( .A0(n16662), .A1(conv_3[343]), .B0(n22615), .B1(conv_3[358]), .Y(n18678) );
  AOI22XL U18583 ( .A0(n36246), .A1(n20553), .B0(n20554), .B1(n22765), .Y(
        n28364) );
  NOR2X1 U18584 ( .A(n27735), .B(n31691), .Y(n23517) );
  NOR2X1 U18585 ( .A(conv_3[410]), .B(n32627), .Y(n19207) );
  AOI22XL U18586 ( .A0(n22369), .A1(n22211), .B0(n22370), .B1(n22204), .Y(
        n19143) );
  NOR2X1 U18587 ( .A(n29426), .B(n31871), .Y(n23066) );
  INVX4 U18588 ( .A(n18777), .Y(n25299) );
  OAI21XL U18589 ( .A0(conv_3[139]), .A1(n23777), .B0(n23776), .Y(n23778) );
  AOI22XL U18590 ( .A0(n19009), .A1(filter_3[23]), .B0(n16676), .B1(
        filter_3[41]), .Y(n18977) );
  NAND2XL U18591 ( .A(n18812), .B(n18811), .Y(n22846) );
  AOI22XL U18592 ( .A0(n34963), .A1(n23244), .B0(n22847), .B1(n23242), .Y(
        n18964) );
  AOI22XL U18593 ( .A0(n19006), .A1(filter_3[6]), .B0(n16676), .B1(
        filter_3[36]), .Y(n19001) );
  NAND4XL U18594 ( .A(n19088), .B(n19087), .C(n19086), .D(n19085), .Y(n23016)
         );
  NAND2XL U18595 ( .A(n18797), .B(n18796), .Y(n22396) );
  NOR2X1 U18596 ( .A(n36199), .B(n36198), .Y(n36200) );
  NOR2X1 U18597 ( .A(affine_2[15]), .B(n36238), .Y(n36199) );
  NOR2X1 U18598 ( .A(affine_2[11]), .B(DP_OP_5170J1_126_4278_n31), .Y(n36169)
         );
  ADDFXL U18599 ( .A(n20632), .B(n20631), .CI(n20630), .CO(n20675), .S(n20671)
         );
  INVXL U18600 ( .A(cursor[6]), .Y(n19182) );
  INVXL U18601 ( .A(n17846), .Y(n17691) );
  NOR2X1 U18602 ( .A(n19182), .B(n16951), .Y(n17444) );
  NOR2X1 U18603 ( .A(n21810), .B(n17172), .Y(n17840) );
  XOR2XL U18604 ( .A(affine_1[24]), .B(n17160), .Y(DP_OP_5166J1_122_9881_n40)
         );
  NAND2XL U18605 ( .A(n26850), .B(n26846), .Y(n20361) );
  NOR2X1 U18606 ( .A(n19703), .B(n17969), .Y(n19709) );
  OAI22XL U18607 ( .A0(n19643), .A1(n19641), .B0(n19640), .B1(n19639), .Y(
        n19729) );
  ADDFXL U18608 ( .A(n28608), .B(n28607), .CI(DP_OP_5171J1_127_4278_n24), .CO(
        n33361), .S(n28613) );
  ADDFXL U18609 ( .A(n28395), .B(n28394), .CI(DP_OP_5170J1_126_4278_n24), .CO(
        n33344), .S(n28400) );
  ADDFXL U18610 ( .A(n28208), .B(n28207), .CI(DP_OP_5169J1_125_4278_n24), .CO(
        n33334), .S(n28213) );
  INVXL U18611 ( .A(n18078), .Y(n19691) );
  INVXL U18612 ( .A(n17929), .Y(n19651) );
  NAND2XL U18613 ( .A(n19242), .B(n19244), .Y(n19632) );
  NOR2X1 U18614 ( .A(ns[2]), .B(ns[1]), .Y(n19243) );
  INVXL U18615 ( .A(n20361), .Y(n36123) );
  NAND4BXL U18616 ( .AN(n18844), .B(n18843), .C(n18842), .D(n18841), .Y(n18845) );
  INVX2 U18617 ( .A(n21730), .Y(n21748) );
  INVX2 U18618 ( .A(n26029), .Y(n26082) );
  NOR2X1 U18619 ( .A(n23462), .B(n23461), .Y(n23463) );
  NOR2X1 U18620 ( .A(n35272), .B(n33524), .Y(n23462) );
  NAND2XL U18621 ( .A(n23587), .B(n24147), .Y(n23969) );
  OR2XL U18622 ( .A(n33403), .B(n25075), .Y(n27031) );
  NOR2XL U18623 ( .A(n30195), .B(n33403), .Y(n27445) );
  INVX2 U18624 ( .A(n21710), .Y(n21764) );
  NOR2X1 U18625 ( .A(n24447), .B(n24446), .Y(n30343) );
  AND2XL U18626 ( .A(n24447), .B(n24446), .Y(n30344) );
  NOR2X1 U18627 ( .A(n35853), .B(n27532), .Y(n30401) );
  AND2X1 U18628 ( .A(n29782), .B(n19109), .Y(n19110) );
  BUFX2 U18629 ( .A(n18912), .Y(n28126) );
  NAND4BXL U18630 ( .AN(n18911), .B(n18910), .C(n18909), .D(n18908), .Y(n18912) );
  AOI22XL U18631 ( .A0(n19009), .A1(filter_2[19]), .B0(n19005), .B1(
        filter_2[13]), .Y(n18909) );
  NOR2X1 U18632 ( .A(n35853), .B(n23793), .Y(n31102) );
  NAND2XL U18633 ( .A(n23579), .B(n24212), .Y(n30406) );
  NOR2X1 U18634 ( .A(n30195), .B(n35853), .Y(n30407) );
  NOR2X1 U18635 ( .A(n27622), .B(n27621), .Y(n30723) );
  NAND2XL U18636 ( .A(n19016), .B(n30789), .Y(n30779) );
  NAND2XL U18637 ( .A(n23604), .B(n30598), .Y(n30622) );
  AOI2BB1XL U18638 ( .A0N(conv_3[316]), .A1N(n30556), .B0(n30557), .Y(n23803)
         );
  NAND2X1 U18639 ( .A(n22110), .B(n30594), .Y(n30574) );
  INVX2 U18640 ( .A(n29680), .Y(n30536) );
  NOR2X1 U18641 ( .A(n34702), .B(n22128), .Y(n22129) );
  NAND2XL U18642 ( .A(n22179), .B(n27496), .Y(n30817) );
  OR2XL U18643 ( .A(n22177), .B(n30536), .Y(n22179) );
  NAND2XL U18644 ( .A(n22907), .B(n27519), .Y(n30793) );
  NAND2XL U18645 ( .A(n22873), .B(n27500), .Y(n30823) );
  BUFX2 U18646 ( .A(n19014), .Y(n29680) );
  NAND4BXL U18647 ( .AN(n19013), .B(n19012), .C(n19011), .D(n19010), .Y(n19014) );
  NOR2X1 U18648 ( .A(n18997), .B(n23203), .Y(n30747) );
  INVX2 U18649 ( .A(n21729), .Y(n21766) );
  NOR2X1 U18650 ( .A(n23640), .B(n23639), .Y(n26939) );
  NOR2X1 U18651 ( .A(n23436), .B(n23435), .Y(n23539) );
  AND2XL U18652 ( .A(n23436), .B(n23435), .Y(n23540) );
  NOR2X1 U18653 ( .A(n23589), .B(n23588), .Y(n23611) );
  AND2XL U18654 ( .A(n23589), .B(n23588), .Y(n23612) );
  AOI2BB1XL U18655 ( .A0N(conv_1[137]), .A1N(n26915), .B0(n26916), .Y(n26748)
         );
  NAND3XL U18656 ( .A(n18832), .B(n18831), .C(n18830), .Y(n18833) );
  OAI2BB2XL U18657 ( .B0(n19227), .B1(n28236), .A0N(n20605), .A1N(filter_1[2]), 
        .Y(n18834) );
  NOR2X1 U18658 ( .A(n22418), .B(n22419), .Y(n26990) );
  AND2XL U18659 ( .A(n22419), .B(n22418), .Y(n26991) );
  AOI2BB1XL U18660 ( .A0N(conv_1[47]), .A1N(n27438), .B0(n27439), .Y(n27326)
         );
  NOR2X1 U18661 ( .A(n26502), .B(n26501), .Y(n27356) );
  AND2XL U18662 ( .A(n26502), .B(n26501), .Y(n27357) );
  NOR2X1 U18663 ( .A(n27738), .B(n27737), .Y(n29547) );
  AND2XL U18664 ( .A(n27738), .B(n27737), .Y(n29548) );
  NOR2X1 U18665 ( .A(n27864), .B(n27863), .Y(n29559) );
  OAI21XL U18666 ( .A0(n29820), .A1(n29815), .B0(n29816), .Y(n28129) );
  NOR2X1 U18667 ( .A(n23076), .B(n23075), .Y(n23991) );
  AND2XL U18668 ( .A(n23076), .B(n23075), .Y(n23992) );
  NAND2XL U18669 ( .A(n23122), .B(n29988), .Y(n23233) );
  NAND2XL U18670 ( .A(n23857), .B(n27411), .Y(n28086) );
  INVX2 U18671 ( .A(n28128), .Y(n35853) );
  NOR2X1 U18672 ( .A(n22970), .B(n22969), .Y(n27851) );
  NAND2X1 U18673 ( .A(n23351), .B(n30413), .Y(n29001) );
  INVXL U18674 ( .A(n25872), .Y(n26081) );
  AND2XL U18675 ( .A(n27624), .B(n27623), .Y(n29632) );
  NOR2X1 U18676 ( .A(n23958), .B(n23957), .Y(n29707) );
  NOR2X1 U18677 ( .A(n23631), .B(n23630), .Y(n29695) );
  AND2XL U18678 ( .A(n23631), .B(n23630), .Y(n29696) );
  NOR2X1 U18679 ( .A(n23606), .B(n23605), .Y(n23766) );
  NAND2XL U18680 ( .A(n30714), .B(n23220), .Y(n23485) );
  NOR2X1 U18681 ( .A(n22144), .B(n22143), .Y(n29689) );
  NOR2X1 U18682 ( .A(n29426), .B(n34426), .Y(n23532) );
  AOI2BB1XL U18683 ( .A0N(conv_3[47]), .A1N(n30747), .B0(n30748), .Y(n29719)
         );
  NOR2X1 U18684 ( .A(n29426), .B(n33988), .Y(n29726) );
  NAND3XL U18685 ( .A(n18994), .B(n18993), .C(n18992), .Y(n18995) );
  OAI2BB1XL U18686 ( .A0N(n20605), .A1N(filter_3[2]), .B0(n18991), .Y(n18996)
         );
  AOI22XL U18687 ( .A0(n19008), .A1(filter_3[44]), .B0(n16676), .B1(
        filter_3[38]), .Y(n18994) );
  NAND2XL U18688 ( .A(n23753), .B(n27509), .Y(n23755) );
  AOI22XL U18689 ( .A0(n25289), .A1(conv_1[64]), .B0(n22690), .B1(conv_1[34]), 
        .Y(n19878) );
  NAND2XL U18690 ( .A(n36246), .B(n22509), .Y(n21535) );
  NAND2X1 U18691 ( .A(n28290), .B(n18204), .Y(n26285) );
  AOI22XL U18692 ( .A0(n34963), .A1(n21543), .B0(n21544), .B1(n24056), .Y(
        n19890) );
  INVX2 U18693 ( .A(n22008), .Y(n21999) );
  AND2XL U18694 ( .A(n23642), .B(n23641), .Y(n27000) );
  NOR2X1 U18695 ( .A(n23642), .B(n23641), .Y(n27001) );
  AND2XL U18696 ( .A(n25252), .B(n25251), .Y(n29571) );
  NOR2X1 U18697 ( .A(n25252), .B(n25251), .Y(n29572) );
  AND2XL U18698 ( .A(n19152), .B(n19151), .Y(n23759) );
  NOR2X1 U18699 ( .A(n19152), .B(n19151), .Y(n23760) );
  AND2XL U18700 ( .A(n22810), .B(n22811), .Y(n30276) );
  NOR2X1 U18701 ( .A(n19216), .B(n19217), .Y(n24224) );
  NOR2X1 U18702 ( .A(n22823), .B(n22824), .Y(n30479) );
  NOR2X1 U18703 ( .A(n22285), .B(n22286), .Y(n30473) );
  AND2XL U18704 ( .A(n23438), .B(n23437), .Y(n24168) );
  NOR2X1 U18705 ( .A(n23438), .B(n23437), .Y(n24169) );
  AND2XL U18706 ( .A(n23591), .B(n23590), .Y(n23975) );
  NOR2X1 U18707 ( .A(n19131), .B(n19130), .Y(n26927) );
  NOR2X1 U18708 ( .A(n24348), .B(n24347), .Y(n32880) );
  AND2XL U18709 ( .A(n25078), .B(n25077), .Y(n27036) );
  NOR2X1 U18710 ( .A(n25078), .B(n25077), .Y(n27037) );
  AOI22XL U18711 ( .A0(n34963), .A1(n25938), .B0(n34961), .B1(n25932), .Y(
        n21867) );
  INVXL U18712 ( .A(n20491), .Y(n22011) );
  OAI222XL U18713 ( .A0(n29021), .A1(n22550), .B0(n22713), .B1(n21858), .C0(
        n19902), .C1(n29033), .Y(n25511) );
  AOI22XL U18714 ( .A0(n25289), .A1(conv_2[394]), .B0(n22690), .B1(conv_2[364]), .Y(n18256) );
  AND2XL U18715 ( .A(n27769), .B(n27768), .Y(n28971) );
  NOR2X1 U18716 ( .A(n27769), .B(n27768), .Y(n28972) );
  NOR2X1 U18717 ( .A(n18934), .B(n18933), .Y(n28989) );
  AND2XL U18718 ( .A(n18934), .B(n18933), .Y(n28990) );
  AND2XL U18719 ( .A(n27740), .B(n27739), .Y(n28983) );
  NOR2X1 U18720 ( .A(n27740), .B(n27739), .Y(n28984) );
  NOR2X1 U18721 ( .A(n27866), .B(n27865), .Y(n28995) );
  OAI21XL U18722 ( .A0(conv_2[408]), .A1(n29420), .B0(n29421), .Y(n28074) );
  AND2XL U18723 ( .A(n23078), .B(n23077), .Y(n29010) );
  NOR2X1 U18724 ( .A(n23124), .B(n23123), .Y(n23356) );
  AND2XL U18725 ( .A(n19113), .B(n19112), .Y(n28870) );
  NOR2X1 U18726 ( .A(n19113), .B(n19112), .Y(n28871) );
  AND2XL U18727 ( .A(n28089), .B(n28090), .Y(n29034) );
  NOR2X1 U18728 ( .A(n28090), .B(n28089), .Y(n29035) );
  NOR2X1 U18729 ( .A(n27853), .B(n27852), .Y(n29040) );
  NOR2X1 U18730 ( .A(n28654), .B(n28653), .Y(n29022) );
  AND2XL U18731 ( .A(n28654), .B(n28653), .Y(n29023) );
  AND2XL U18732 ( .A(n29005), .B(n29004), .Y(n29833) );
  NOR2X1 U18733 ( .A(n29004), .B(n29005), .Y(n29832) );
  NOR2X1 U18734 ( .A(n23480), .B(n23479), .Y(n28741) );
  AND2XL U18735 ( .A(n23480), .B(n23479), .Y(n28740) );
  NOR2X1 U18736 ( .A(n27706), .B(n27705), .Y(n29702) );
  NOR2X1 U18737 ( .A(n24827), .B(n25123), .Y(n18493) );
  NOR2X1 U18738 ( .A(n35107), .B(n25123), .Y(n18499) );
  AOI211XL U18739 ( .A0(n34963), .A1(n35101), .B0(n28306), .C0(n28305), .Y(
        n28308) );
  NAND2X1 U18740 ( .A(n26470), .B(n36245), .Y(n35196) );
  NOR2X1 U18741 ( .A(n23960), .B(n23959), .Y(n31926) );
  AND2XL U18742 ( .A(n23960), .B(n23959), .Y(n31925) );
  AND2XL U18743 ( .A(n23633), .B(n23632), .Y(n32019) );
  NOR2X1 U18744 ( .A(n23633), .B(n23632), .Y(n32018) );
  AND2XL U18745 ( .A(n23509), .B(n23508), .Y(n31626) );
  NOR2X1 U18746 ( .A(n23509), .B(n23508), .Y(n31625) );
  OAI21XL U18747 ( .A0(conv_3[333]), .A1(n23766), .B0(n23765), .Y(n23767) );
  OR2XL U18748 ( .A(n23805), .B(n23804), .Y(n23811) );
  NOR2X1 U18749 ( .A(n22861), .B(n22860), .Y(n26328) );
  AND2XL U18750 ( .A(n22133), .B(n22132), .Y(n26316) );
  NOR2X1 U18751 ( .A(n22133), .B(n22132), .Y(n26315) );
  NOR2X1 U18752 ( .A(n31691), .B(n22257), .Y(n29070) );
  NOR2X1 U18753 ( .A(n22183), .B(n22182), .Y(n29746) );
  AND2XL U18754 ( .A(n22183), .B(n22182), .Y(n29745) );
  NOR2X1 U18755 ( .A(n23534), .B(n23533), .Y(n23777) );
  AND2XL U18756 ( .A(n23690), .B(n23689), .Y(n28950) );
  NOR2X1 U18757 ( .A(n23690), .B(n23689), .Y(n28949) );
  OAI21XL U18758 ( .A0(conv_3[108]), .A1(n29650), .B0(n29651), .Y(n22910) );
  AOI2BB1XL U18759 ( .A0N(conv_1[534]), .A1N(n29214), .B0(n29236), .Y(n29189)
         );
  INVX3 U18760 ( .A(n22765), .Y(n36246) );
  INVXL U18761 ( .A(n28418), .Y(n26632) );
  AOI22XL U18762 ( .A0(n28528), .A1(n28412), .B0(n34963), .B1(n28410), .Y(
        n25314) );
  NOR4BXL U18763 ( .AN(n25429), .B(n25428), .C(n25427), .D(n25426), .Y(n25430)
         );
  INVX2 U18764 ( .A(n19401), .Y(n21011) );
  NOR2X1 U18765 ( .A(conv_1[518]), .B(n27257), .Y(n25262) );
  AND2XL U18766 ( .A(n30267), .B(n24912), .Y(n27260) );
  NAND4XL U18767 ( .A(n18865), .B(n18864), .C(n18863), .D(n18862), .Y(n22151)
         );
  NAND4XL U18768 ( .A(n18877), .B(n18876), .C(n18875), .D(n18874), .Y(n22152)
         );
  NOR2X1 U18769 ( .A(n30325), .B(n35534), .Y(n30326) );
  NOR2X1 U18770 ( .A(conv_1[491]), .B(n30324), .Y(n30325) );
  AOI2BB1XL U18771 ( .A0N(conv_1[487]), .A1N(n35532), .B0(n35534), .Y(n35539)
         );
  NOR2X1 U18772 ( .A(n35536), .B(n35533), .Y(n35540) );
  AOI2BB1XL U18773 ( .A0N(conv_1[469]), .A1N(n27006), .B0(n27007), .Y(n18855)
         );
  NOR2X1 U18774 ( .A(conv_1[459]), .B(n30031), .Y(n27239) );
  AOI2BB1XL U18775 ( .A0N(conv_1[440]), .A1N(n27166), .B0(n27149), .Y(n27154)
         );
  NOR2X1 U18776 ( .A(n27167), .B(n27171), .Y(n27155) );
  NOR2X1 U18777 ( .A(n33393), .B(n29328), .Y(n29221) );
  AOI2BB1XL U18778 ( .A0N(conv_1[379]), .A1N(n23759), .B0(n23760), .Y(n19153)
         );
  NOR2X1 U18779 ( .A(n25274), .B(n25270), .Y(n29385) );
  NOR2X1 U18780 ( .A(conv_1[307]), .B(n19218), .Y(n22318) );
  AOI2BB1XL U18781 ( .A0N(conv_1[294]), .A1N(n23182), .B0(n22827), .Y(n23187)
         );
  AOI2BB1XL U18782 ( .A0N(conv_1[291]), .A1N(n29376), .B0(n22827), .Y(n23170)
         );
  AOI2BB1XL U18783 ( .A0N(conv_1[290]), .A1N(n29311), .B0(n22827), .Y(n29376)
         );
  NOR2X1 U18784 ( .A(n29310), .B(n29315), .Y(n29377) );
  NAND2XL U18785 ( .A(n27632), .B(n34455), .Y(n22827) );
  AOI2BB1XL U18786 ( .A0N(conv_1[276]), .A1N(n29316), .B0(n29339), .Y(n29344)
         );
  NOR2X1 U18787 ( .A(n29317), .B(n29321), .Y(n29345) );
  NOR2X1 U18788 ( .A(n29339), .B(n22287), .Y(n29370) );
  AOI2BB1XL U18789 ( .A0N(conv_1[234]), .A1N(n35405), .B0(n34276), .Y(n31127)
         );
  NOR2X1 U18790 ( .A(n35403), .B(n35407), .Y(n31128) );
  AOI2BB1XL U18791 ( .A0N(conv_1[229]), .A1N(n23909), .B0(n23910), .Y(n22299)
         );
  AOI2BB1XL U18792 ( .A0N(conv_1[187]), .A1N(n23599), .B0(n32988), .Y(n35357)
         );
  NOR2X1 U18793 ( .A(n23598), .B(n23597), .Y(n35358) );
  AOI2BB1XL U18794 ( .A0N(conv_1[184]), .A1N(n23975), .B0(n23976), .Y(n23593)
         );
  NOR2X1 U18795 ( .A(n27540), .B(n27538), .Y(n23935) );
  AOI2BB1XL U18796 ( .A0N(n23404), .A1N(n23400), .B0(n34044), .Y(n23406) );
  AOI2BB1XL U18797 ( .A0N(conv_1[155]), .A1N(n23399), .B0(n23394), .Y(n23405)
         );
  AOI2BB1XL U18798 ( .A0N(conv_1[139]), .A1N(n26927), .B0(n26928), .Y(n19132)
         );
  NAND2XL U18799 ( .A(n18805), .B(n18804), .Y(n22844) );
  AOI2BB1XL U18800 ( .A0N(conv_1[95]), .A1N(n26779), .B0(n31334), .Y(n26789)
         );
  AOI2BB1XL U18801 ( .A0N(conv_1[85]), .A1N(n26724), .B0(n26735), .Y(n26729)
         );
  OAI2BB1XL U18802 ( .A0N(n35316), .A1N(conv_1[50]), .B0(n26132), .Y(n26134)
         );
  AOI2BB1XL U18803 ( .A0N(conv_1[49]), .A1N(n27456), .B0(n27457), .Y(n26133)
         );
  NOR2X1 U18804 ( .A(n30587), .B(n30588), .Y(n30589) );
  NOR2X1 U18805 ( .A(n33372), .B(n29095), .Y(n29101) );
  INVXL U18806 ( .A(n16672), .Y(n28559) );
  NOR2X1 U18807 ( .A(n26575), .B(n20726), .Y(n21765) );
  OR2X1 U18808 ( .A(n16721), .B(n20726), .Y(n22018) );
  OR4XL U18809 ( .A(n26100), .B(n26099), .C(n26098), .D(n26097), .Y(n26107) );
  AOI22XL U18810 ( .A0(n25306), .A1(conv_2[285]), .B0(n16673), .B1(conv_2[315]), .Y(n20730) );
  AOI22XL U18811 ( .A0(n25306), .A1(conv_2[105]), .B0(n16673), .B1(conv_2[135]), .Y(n20728) );
  AOI22XL U18812 ( .A0(n25306), .A1(conv_2[45]), .B0(n16662), .B1(conv_2[60]), 
        .Y(n20738) );
  AOI22XL U18813 ( .A0(n25306), .A1(conv_2[165]), .B0(n16662), .B1(conv_2[180]), .Y(n20736) );
  OR2XL U18814 ( .A(n36245), .B(n35241), .Y(n26474) );
  BUFX2 U18815 ( .A(n16702), .Y(n26374) );
  OR2XL U18816 ( .A(N18471), .B(n18205), .Y(n35200) );
  AND2XL U18817 ( .A(n36088), .B(n18935), .Y(n31017) );
  NOR2X1 U18818 ( .A(n36088), .B(n18935), .Y(n31016) );
  NOR2X1 U18819 ( .A(n33601), .B(n34130), .Y(n27758) );
  AOI21XL U18820 ( .A0(n33602), .A1(conv_2[486]), .B0(n34132), .Y(n27759) );
  NOR2X1 U18821 ( .A(conv_2[471]), .B(n27872), .Y(n27874) );
  AOI2BB1XL U18822 ( .A0N(conv_2[442]), .A1N(n28935), .B0(n28937), .Y(n36065)
         );
  AOI2BB1XL U18823 ( .A0N(conv_2[411]), .A1N(n29486), .B0(n33321), .Y(n28082)
         );
  NOR2X1 U18824 ( .A(n29487), .B(n29491), .Y(n28081) );
  OAI21XL U18825 ( .A0(conv_2[409]), .A1(n28858), .B0(n28859), .Y(n28076) );
  INVXL U18826 ( .A(n34634), .Y(n33953) );
  NOR2X1 U18827 ( .A(n35997), .B(n23086), .Y(n28096) );
  AOI21XL U18828 ( .A0(n28058), .A1(n28057), .B0(n33079), .Y(n28063) );
  NOR2X1 U18829 ( .A(n28058), .B(n28056), .Y(n28064) );
  NOR2X1 U18830 ( .A(n35981), .B(n35985), .Y(n28045) );
  NOR2X1 U18831 ( .A(n35969), .B(n35972), .Y(n28627) );
  AOI2BB1XL U18832 ( .A0N(conv_2[307]), .A1N(n28898), .B0(n35970), .Y(n29946)
         );
  AOI2BB1XL U18833 ( .A0N(conv_2[305]), .A1N(n30857), .B0(n35970), .Y(n28917)
         );
  NOR2X1 U18834 ( .A(n30858), .B(n30861), .Y(n28918) );
  AOI2BB1XL U18835 ( .A0N(conv_2[291]), .A1N(n35955), .B0(n33135), .Y(n30917)
         );
  OAI211XL U18836 ( .A0(n21095), .A1(n19181), .B0(n19140), .C0(n19139), .Y(
        n22850) );
  AOI22XL U18837 ( .A0(n22369), .A1(n22397), .B0(n21100), .B1(n22212), .Y(
        n19140) );
  INVXL U18838 ( .A(n35957), .Y(n33135) );
  NOR2X1 U18839 ( .A(conv_2[261]), .B(n34599), .Y(n19044) );
  AOI2BB1XL U18840 ( .A0N(conv_2[246]), .A1N(n29143), .B0(n29455), .Y(n29167)
         );
  NOR2X1 U18841 ( .A(n29148), .B(n29144), .Y(n29168) );
  OAI21XL U18842 ( .A0(conv_2[244]), .A1(n28977), .B0(n28978), .Y(n28149) );
  NOR2X1 U18843 ( .A(n29862), .B(n29867), .Y(n29857) );
  AOI2BB1XL U18844 ( .A0N(conv_2[140]), .A1N(n34240), .B0(n35899), .Y(n30076)
         );
  NOR2X1 U18845 ( .A(n30136), .B(n30135), .Y(n30149) );
  AND2XL U18846 ( .A(n30204), .B(n30944), .Y(n30205) );
  AOI222XL U18847 ( .A0(n24015), .A1(n24016), .B0(n24015), .B1(conv_2[94]), 
        .C0(n24016), .C1(conv_2[94]), .Y(n19171) );
  AOI2BB1XL U18848 ( .A0N(conv_2[70]), .A1N(n30125), .B0(n30242), .Y(n30240)
         );
  NOR2X1 U18849 ( .A(n28715), .B(n28714), .Y(n27826) );
  NOR2X1 U18850 ( .A(n27716), .B(n27712), .Y(n27718) );
  AOI2BB1XL U18851 ( .A0N(conv_2[37]), .A1N(n27711), .B0(n35862), .Y(n27717)
         );
  AOI2BB1XL U18852 ( .A0N(conv_2[34]), .A1N(n29701), .B0(n29702), .Y(n27707)
         );
  NAND4BX1 U18853 ( .AN(n18918), .B(n18917), .C(n18916), .D(n18915), .Y(n28124) );
  AOI22XL U18854 ( .A0(n19009), .A1(filter_2[18]), .B0(n19006), .B1(
        filter_2[6]), .Y(n18916) );
  AOI22XL U18855 ( .A0(n19008), .A1(filter_2[42]), .B0(n19004), .B1(
        filter_2[30]), .Y(n18915) );
  OAI2BB1XL U18856 ( .A0N(counter[3]), .A1N(filter_2[48]), .B0(n18914), .Y(
        n18918) );
  AOI2BB1XL U18857 ( .A0N(conv_2[19]), .A1N(n29713), .B0(n29714), .Y(n27555)
         );
  NOR2X1 U18858 ( .A(n28957), .B(n28959), .Y(n31141) );
  NOR2X1 U18859 ( .A(n28961), .B(n28960), .Y(n31142) );
  INVXL U18860 ( .A(n21536), .Y(n21763) );
  INVXL U18861 ( .A(n21237), .Y(n21761) );
  AOI211XL U18862 ( .A0(n34963), .A1(n21432), .B0(n20565), .C0(n20564), .Y(
        n20570) );
  NOR2X1 U18863 ( .A(n20538), .B(n21960), .Y(n20540) );
  AOI22XL U18864 ( .A0(n25289), .A1(conv_3[180]), .B0(n22690), .B1(conv_3[150]), .Y(n19262) );
  INVXL U18865 ( .A(n22009), .Y(n34952) );
  INVXL U18866 ( .A(n22018), .Y(n21992) );
  AOI22XL U18867 ( .A0(n34963), .A1(n35168), .B0(n35169), .B1(n26451), .Y(
        n24816) );
  NOR4BBXL U18868 ( .AN(n24898), .BN(n24897), .C(n24896), .D(n24895), .Y(
        n24899) );
  INVXL U18869 ( .A(n28391), .Y(n35229) );
  NOR2X2 U18870 ( .A(n26479), .B(n25123), .Y(n18463) );
  NOR2X1 U18871 ( .A(n32065), .B(n33918), .Y(n32082) );
  NOR2X1 U18872 ( .A(n32064), .B(n32063), .Y(n32083) );
  NOR2X1 U18873 ( .A(n33759), .B(n35789), .Y(n31950) );
  AOI2BB1XL U18874 ( .A0N(conv_3[440]), .A1N(n31933), .B0(n35789), .Y(n31938)
         );
  INVX2 U18875 ( .A(n18757), .Y(n21100) );
  INVXL U18876 ( .A(n28407), .Y(n18757) );
  AOI22XL U18877 ( .A0(n22369), .A1(n19052), .B0(n22370), .B1(n19051), .Y(
        n23252) );
  NOR2X1 U18878 ( .A(conv_3[416]), .B(n32011), .Y(n31994) );
  NOR2X1 U18879 ( .A(n19207), .B(n32558), .Y(n32004) );
  NOR2X1 U18880 ( .A(n19207), .B(n32626), .Y(n32005) );
  NOR2X1 U18881 ( .A(conv_3[401]), .B(n33220), .Y(n33222) );
  AOI2BB1XL U18882 ( .A0N(conv_3[396]), .A1N(n32032), .B0(n33695), .Y(n32038)
         );
  AOI2BB1XL U18883 ( .A0N(conv_3[395]), .A1N(n32026), .B0(n33695), .Y(n32032)
         );
  AOI2BB1XL U18884 ( .A0N(conv_3[385]), .A1N(n31461), .B0(n32200), .Y(n32197)
         );
  AOI2BB1XL U18885 ( .A0N(conv_3[367]), .A1N(n31654), .B0(n35761), .Y(n31648)
         );
  AOI2BB1XL U18886 ( .A0N(conv_3[365]), .A1N(n31637), .B0(n35761), .Y(n31660)
         );
  NOR2X1 U18887 ( .A(n31636), .B(n31641), .Y(n31661) );
  AOI2BB1XL U18888 ( .A0N(conv_3[350]), .A1N(n31480), .B0(n32130), .Y(n31450)
         );
  NOR2X1 U18889 ( .A(n31479), .B(n31484), .Y(n31449) );
  NOR2X1 U18890 ( .A(n31957), .B(n31956), .Y(n31975) );
  OAI21XL U18891 ( .A0(conv_3[334]), .A1(n26945), .B0(n26946), .Y(n23769) );
  AOI2BB1XL U18892 ( .A0N(conv_3[325]), .A1N(n31915), .B0(n33281), .Y(n31919)
         );
  AOI222XL U18893 ( .A0(n28756), .A1(conv_3[319]), .B0(n28756), .B1(n28755), 
        .C0(conv_3[319]), .C1(n28755), .Y(n28757) );
  NOR2X1 U18894 ( .A(n35731), .B(n35735), .Y(n31496) );
  AOI2BB1XL U18895 ( .A0N(conv_3[280]), .A1N(n31757), .B0(n32599), .Y(n31762)
         );
  NOR2X1 U18896 ( .A(n35648), .B(n31848), .Y(n31865) );
  NOR2X1 U18897 ( .A(conv_3[176]), .B(n31577), .Y(n31579) );
  AOI2BB1XL U18898 ( .A0N(conv_3[175]), .A1N(n35637), .B0(n32221), .Y(n31577)
         );
  NOR2X1 U18899 ( .A(conv_3[159]), .B(n32297), .Y(n32251) );
  AOI2BB1XL U18900 ( .A0N(conv_3[158]), .A1N(n32278), .B0(n32252), .Y(n32297)
         );
  NOR2X1 U18901 ( .A(n32248), .B(n32252), .Y(n32278) );
  NOR2X1 U18902 ( .A(n32250), .B(n32249), .Y(n32279) );
  NAND4X1 U18903 ( .A(n18889), .B(n18888), .C(n18887), .D(n18886), .Y(n22153)
         );
  AOI22XL U18904 ( .A0(pixel[24]), .A1(n19099), .B0(pixel[20]), .B1(n16734), 
        .Y(n18887) );
  AOI22XL U18905 ( .A0(pixel[22]), .A1(n21887), .B0(pixel[26]), .B1(n19098), 
        .Y(n18886) );
  AOI22XL U18906 ( .A0(pixel[23]), .A1(n19475), .B0(pixel[25]), .B1(n19097), 
        .Y(n18889) );
  NAND4XL U18907 ( .A(n18869), .B(n18868), .C(n18867), .D(n18866), .Y(n22266)
         );
  AOI2BB1XL U18908 ( .A0N(conv_3[112]), .A1N(n31797), .B0(n31786), .Y(n31791)
         );
  AOI21XL U18909 ( .A0(n31798), .A1(conv_3[112]), .B0(n34196), .Y(n31792) );
  OAI21XL U18910 ( .A0(conv_3[109]), .A1(n31768), .B0(n31767), .Y(n31769) );
  AOI2BB1XL U18911 ( .A0N(conv_3[97]), .A1N(n31673), .B0(n35615), .Y(n31685)
         );
  NOR2X1 U18912 ( .A(n31678), .B(n31674), .Y(n31686) );
  AOI2BB1XL U18913 ( .A0N(conv_3[82]), .A1N(n31833), .B0(n35607), .Y(n31810)
         );
  NOR2X1 U18914 ( .A(n31838), .B(n31834), .Y(n31811) );
  AOI2BB1XL U18915 ( .A0N(conv_3[80]), .A1N(n34151), .B0(n35607), .Y(n31821)
         );
  NOR2X1 U18916 ( .A(n34150), .B(n34154), .Y(n31822) );
  NAND2XL U18917 ( .A(n19031), .B(n19030), .Y(n22403) );
  AOI22XL U18918 ( .A0(n35181), .A1(n22846), .B0(n28556), .B1(n22845), .Y(
        n22406) );
  NAND2XL U18919 ( .A(n18799), .B(n18798), .Y(n22402) );
  NAND2XL U18920 ( .A(n19029), .B(n19028), .Y(n23089) );
  AOI22XL U18921 ( .A0(n22370), .A1(n22210), .B0(n21100), .B1(n22211), .Y(
        n19029) );
  AOI22XL U18922 ( .A0(n22362), .A1(n22212), .B0(n22369), .B1(n22889), .Y(
        n19028) );
  NOR2X1 U18923 ( .A(conv_3[56]), .B(n32176), .Y(n32179) );
  AOI2BB1XL U18924 ( .A0N(conv_3[55]), .A1N(n31216), .B0(n32178), .Y(n32176)
         );
  AOI2BB1XL U18925 ( .A0N(conv_3[51]), .A1N(n31211), .B0(n32178), .Y(n31204)
         );
  NAND4XL U18926 ( .A(n18881), .B(n18880), .C(n18879), .D(n18878), .Y(n22448)
         );
  AOI22XL U18927 ( .A0(pixel[37]), .A1(n22021), .B0(pixel[42]), .B1(n19098), 
        .Y(n18880) );
  NAND4XL U18928 ( .A(n18873), .B(n18872), .C(n18871), .D(n18870), .Y(n22447)
         );
  AOI22XL U18929 ( .A0(n23272), .A1(n22266), .B0(n23274), .B1(n22151), .Y(
        n22155) );
  AOI22XL U18930 ( .A0(n23278), .A1(n22153), .B0(n23276), .B1(n22152), .Y(
        n22154) );
  NAND4XL U18931 ( .A(n18893), .B(n18892), .C(n18891), .D(n18890), .Y(n22449)
         );
  NAND4XL U18932 ( .A(n18885), .B(n18884), .C(n18883), .D(n18882), .Y(n22450)
         );
  INVXL U18933 ( .A(n33824), .Y(n32178) );
  OAI21XL U18934 ( .A0(conv_3[34]), .A1(n29663), .B0(n29664), .Y(n24470) );
  NAND4XL U18935 ( .A(n19103), .B(n19102), .C(n19101), .D(n19100), .Y(n23784)
         );
  NAND4XL U18936 ( .A(n19084), .B(n19083), .C(n19082), .D(n19081), .Y(n23781)
         );
  NAND4XL U18937 ( .A(n19076), .B(n19075), .C(n19074), .D(n19073), .Y(n23782)
         );
  AOI22XL U18938 ( .A0(pixel[42]), .A1(n21954), .B0(pixel[45]), .B1(n21887), 
        .Y(n19073) );
  OAI211XL U18939 ( .A0(n23282), .A1(n23281), .B0(n23280), .C0(n23279), .Y(
        n23786) );
  NOR2X1 U18940 ( .A(n20363), .B(n20362), .Y(n30349) );
  NAND2X1 U18941 ( .A(n36244), .B(n16700), .Y(n23052) );
  AND2XL U18942 ( .A(counter[6]), .B(counter[5]), .Y(n26850) );
  NAND2XL U18943 ( .A(counter[3]), .B(counter[4]), .Y(n20164) );
  NAND3BXL U18944 ( .AN(n18186), .B(cs[0]), .C(n18185), .Y(n18188) );
  NAND2XL U18945 ( .A(cs[1]), .B(cs[2]), .Y(n18186) );
  INVXL U18946 ( .A(n20165), .Y(n18158) );
  NAND2XL U18947 ( .A(counter[2]), .B(n19229), .Y(n18172) );
  ADDFXL U18948 ( .A(DP_OP_5168J1_124_9881_n16), .B(DP_OP_5168J1_124_9881_n14), 
        .CI(n33069), .CO(n33070), .S(n22251) );
  ADDFXL U18949 ( .A(DP_OP_5168J1_124_9881_n21), .B(DP_OP_5168J1_124_9881_n17), 
        .CI(n22249), .CO(n33069), .S(n21093) );
  OAI21XL U18950 ( .A0(affine_1[9]), .A1(n20638), .B0(n33075), .Y(n22250) );
  OAI21XL U18951 ( .A0(affine_1[19]), .A1(n20638), .B0(n33075), .Y(n25243) );
  ADDFXL U18952 ( .A(n20700), .B(n20699), .CI(n20698), .CO(n20678), .S(n20701)
         );
  OAI21XL U18953 ( .A0(affine_1[29]), .A1(n20638), .B0(n33075), .Y(n25069) );
  NOR2X1 U18954 ( .A(n20616), .B(n20615), .Y(n33563) );
  NOR3X1 U18955 ( .A(n20600), .B(n20361), .C(n20599), .Y(n36155) );
  INVXL U18956 ( .A(n36155), .Y(n36153) );
  INVXL U18957 ( .A(n16647), .Y(n32967) );
  NAND2XL U18958 ( .A(counter[4]), .B(n26850), .Y(n26851) );
  AOI21X1 U18959 ( .A0(n26849), .A1(n26848), .B0(n26847), .Y(n26852) );
  AND2X1 U18960 ( .A(n20360), .B(n20359), .Y(n20419) );
  NOR3XL U18961 ( .A(n20358), .B(n20362), .C(n20361), .Y(n20359) );
  ADDFXL U18962 ( .A(n33361), .B(n33360), .CI(n33359), .CO(n33362), .S(n28614)
         );
  NAND2XL U18963 ( .A(weight_2_bias_1[5]), .B(n20614), .Y(n33368) );
  ADDFXL U18964 ( .A(n33334), .B(n33333), .CI(n33332), .CO(n33335), .S(n28214)
         );
  ADDFXL U18965 ( .A(DP_OP_5169J1_125_4278_n26), .B(DP_OP_5169J1_125_4278_n28), 
        .CI(n24547), .CO(n28212), .S(n20719) );
  ADDFXL U18966 ( .A(DP_OP_5169J1_125_4278_n33), .B(DP_OP_5169J1_125_4278_n29), 
        .CI(n20718), .CO(n24547), .S(n20356) );
  ADDFXL U18967 ( .A(DP_OP_5169J1_125_4278_n34), .B(DP_OP_5169J1_125_4278_n38), 
        .CI(n20355), .CO(n20718), .S(n20148) );
  NAND2XL U18968 ( .A(weight_2_bias_3[5]), .B(n20614), .Y(n33340) );
  NAND2X1 U18969 ( .A(n36123), .B(n36122), .Y(n36136) );
  NOR4XL U18970 ( .A(counter[4]), .B(n20605), .C(n20604), .D(n30350), .Y(
        n20608) );
  NOR4XL U18971 ( .A(n21514), .B(n21513), .C(n21512), .D(n21511), .Y(n34812)
         );
  AOI211XL U18972 ( .A0(n28465), .A1(n20218), .B0(n19852), .C0(n19851), .Y(
        n34797) );
  AOI211XL U18973 ( .A0(n34992), .A1(n26546), .B0(n25406), .C0(n25405), .Y(
        n34790) );
  AOI22XL U18974 ( .A0(n26263), .A1(n26395), .B0(n34963), .B1(n25392), .Y(
        n25404) );
  AOI211XL U18975 ( .A0(n34992), .A1(n26547), .B0(n26397), .C0(n26396), .Y(
        n34803) );
  AOI21XL U18976 ( .A0(n26391), .A1(n26390), .B0(N18014), .Y(n26397) );
  AOI211XL U18977 ( .A0(n34827), .A1(n26554), .B0(n26553), .C0(n26552), .Y(
        n34807) );
  NOR2XL U18978 ( .A(n26550), .B(n35159), .Y(n24629) );
  NOR4BXL U18979 ( .AN(n22700), .B(n22699), .C(n22698), .D(n22697), .Y(n34836)
         );
  OAI22XL U18980 ( .A0(n27232), .A1(n27644), .B0(n27421), .B1(n27429), .Y(
        n27435) );
  NOR2X1 U18981 ( .A(n35272), .B(n30648), .Y(n30666) );
  AOI211XL U18982 ( .A0(n35272), .A1(n22291), .B0(n22290), .C0(n29136), .Y(
        n23951) );
  OAI32XL U18983 ( .A0(n23433), .A1(n27848), .A2(n35272), .B0(n27429), .B1(
        n24216), .Y(n24221) );
  OAI22XL U18984 ( .A0(n23586), .A1(n34703), .B0(n24137), .B1(n27429), .Y(
        n24148) );
  OAI22XL U18985 ( .A0(n26499), .A1(n30195), .B0(n27429), .B1(n26498), .Y(
        n27463) );
  NAND2X1 U18986 ( .A(n22896), .B(filter_1_bias[1]), .Y(n33067) );
  NOR4BXL U18987 ( .AN(n21025), .B(n21024), .C(n21023), .D(n21022), .Y(n34887)
         );
  AOI211XL U18988 ( .A0(n16755), .A1(n25889), .B0(n25888), .C0(n25887), .Y(
        n26113) );
  AOI211XL U18989 ( .A0(n28465), .A1(n25889), .B0(n21855), .C0(n21854), .Y(
        n34868) );
  AOI211XL U18990 ( .A0(n26263), .A1(n25115), .B0(n24975), .C0(n24974), .Y(
        n34863) );
  AOI22XL U18991 ( .A0(n16667), .A1(n25114), .B0(n34963), .B1(n24972), .Y(
        n24973) );
  AOI211XL U18992 ( .A0(n24714), .A1(n26470), .B0(n24713), .C0(n24712), .Y(
        n34881) );
  AOI22XL U18993 ( .A0(n34963), .A1(n25115), .B0(n16670), .B1(n25114), .Y(
        n24710) );
  AOI211XL U18994 ( .A0(n16755), .A1(n24714), .B0(n18397), .C0(n18396), .Y(
        n22200) );
  AOI211XL U18995 ( .A0(n28324), .A1(n25487), .B0(n25486), .C0(n25485), .Y(
        n34898) );
  NAND2XL U18996 ( .A(n30299), .B(conv_2[376]), .Y(n30298) );
  AOI221XL U18997 ( .A0(n18913), .A1(n23853), .B0(n28126), .B1(n34453), .C0(
        n31871), .Y(n30303) );
  NOR2X1 U18998 ( .A(n18913), .B(n29768), .Y(n29770) );
  OAI32XL U18999 ( .A0(n34431), .A1(n22257), .A2(n18913), .B0(n28126), .B1(
        n23347), .Y(n31091) );
  NOR2X1 U19000 ( .A(n18913), .B(n23574), .Y(n23229) );
  NOR2X1 U19001 ( .A(conv_2[61]), .B(n35844), .Y(n35850) );
  NOR2X1 U19002 ( .A(n24268), .B(n24270), .Y(n24266) );
  NAND2X1 U19003 ( .A(n22896), .B(filter_2_bias[1]), .Y(n35847) );
  NOR4XL U19004 ( .A(n21166), .B(n21165), .C(n21164), .D(n21163), .Y(n35011)
         );
  AOI211XL U19005 ( .A0(n16755), .A1(n20451), .B0(n19517), .C0(n19516), .Y(
        n35023) );
  AOI211XL U19006 ( .A0(n28465), .A1(n20451), .B0(n20450), .C0(n20449), .Y(
        n34975) );
  OAI2BB1XL U19007 ( .A0N(n34963), .A1N(n26179), .B0(n26178), .Y(n26180) );
  AOI22XL U19008 ( .A0(n16659), .A1(n35154), .B0(n34963), .B1(n35152), .Y(
        n24846) );
  OAI211XL U19009 ( .A0(n28301), .A1(n28304), .B0(n28300), .C0(n28299), .Y(
        n35004) );
  AOI211XL U19010 ( .A0(n34963), .A1(n35151), .B0(n28298), .C0(n28297), .Y(
        n28299) );
  NOR2X1 U19011 ( .A(n35157), .B(n28349), .Y(n28298) );
  AOI211XL U19012 ( .A0(n16664), .A1(n25715), .B0(n25714), .C0(n25713), .Y(
        n26702) );
  NOR2X1 U19013 ( .A(n35157), .B(n26621), .Y(n25714) );
  OAI32XL U19014 ( .A0(n19015), .A1(n27860), .A2(n30536), .B0(n29680), .B1(
        n31376), .Y(n30790) );
  AOI211XL U19015 ( .A0(n30536), .A1(n23216), .B0(n23215), .C0(n19108), .Y(
        n31023) );
  OAI32XL U19016 ( .A0(n22109), .A1(n28721), .A2(n30536), .B0(n29680), .B1(
        n30606), .Y(n30595) );
  OAI22XL U19017 ( .A0(n22178), .A1(n23296), .B0(n22177), .B1(n29680), .Y(
        n27497) );
  OAI32XL U19018 ( .A0(n22906), .A1(n34715), .A2(n30536), .B0(n29680), .B1(
        n30829), .Y(n27520) );
  OAI22XL U19019 ( .A0(n22872), .A1(n26509), .B0(n29680), .B1(n30833), .Y(
        n27501) );
  NAND2XL U19020 ( .A(n29680), .B(n30833), .Y(n22872) );
  NOR2X1 U19021 ( .A(n21110), .B(n21108), .Y(n29428) );
  NAND2X1 U19022 ( .A(n22896), .B(filter_3_bias[1]), .Y(n33550) );
  NAND4XL U19023 ( .A(n20234), .B(n20233), .C(n20232), .D(n20231), .Y(n34842)
         );
  OAI2BB1XL U19024 ( .A0N(n16700), .A1N(n20230), .B0(n19829), .Y(n34799) );
  AOI211XL U19025 ( .A0(n34954), .A1(n21520), .B0(n19828), .C0(n19827), .Y(
        n19829) );
  OAI211XL U19026 ( .A0(n26555), .A1(n34958), .B0(n25391), .C0(n25390), .Y(
        n34792) );
  AOI211XL U19027 ( .A0(n34963), .A1(n26398), .B0(n25389), .C0(n25388), .Y(
        n25391) );
  OAI211XL U19028 ( .A0(n34989), .A1(n26557), .B0(n26405), .C0(n26404), .Y(
        n34804) );
  AOI22XL U19029 ( .A0(n34963), .A1(n26399), .B0(n16670), .B1(n26398), .Y(
        n26405) );
  AOI211XL U19030 ( .A0(n26562), .A1(n26451), .B0(n26403), .C0(n26402), .Y(
        n26404) );
  AOI211XL U19031 ( .A0(n26562), .A1(n26561), .B0(n26560), .C0(n26559), .Y(
        n26565) );
  NAND2XL U19032 ( .A(n27233), .B(n27434), .Y(n27379) );
  OR2XL U19033 ( .A(n27421), .B(n35272), .Y(n27233) );
  NOR2X1 U19034 ( .A(n23724), .B(n23723), .Y(n23726) );
  NOR2X1 U19035 ( .A(n33403), .B(n29761), .Y(n29763) );
  ADDFXL U19036 ( .A(conv_1[332]), .B(n22980), .CI(n22979), .CO(n22981), .S(
        n22943) );
  NOR2X1 U19037 ( .A(n30480), .B(n30479), .Y(n30482) );
  NOR2X1 U19038 ( .A(n30474), .B(n30473), .Y(n30476) );
  NOR2X1 U19039 ( .A(n26916), .B(n26915), .Y(n26918) );
  NOR2X1 U19040 ( .A(n33403), .B(n30466), .Y(n30468) );
  NOR2X1 U19041 ( .A(n26685), .B(n26684), .Y(n26687) );
  NOR2X1 U19042 ( .A(n26991), .B(n26990), .Y(n26993) );
  NOR2X1 U19043 ( .A(n27439), .B(n27438), .Y(n27441) );
  NOR2XL U19044 ( .A(n33403), .B(n35857), .Y(intadd_2_B_0_) );
  NAND2X1 U19045 ( .A(n22896), .B(filter_1_bias[2]), .Y(n33542) );
  OAI2BB1XL U19046 ( .A0N(n16755), .A1N(n25869), .B0(n25868), .Y(n34924) );
  AOI211XL U19047 ( .A0(n26081), .A1(n25867), .B0(n25866), .C0(n25865), .Y(
        n25868) );
  OAI2BB1XL U19048 ( .A0N(n16700), .A1N(n25869), .B0(n21840), .Y(n34869) );
  AOI211XL U19049 ( .A0(n16667), .A1(n25859), .B0(n21839), .C0(n21838), .Y(
        n21840) );
  OAI21XL U19050 ( .A0(n25128), .A1(n28467), .B0(n24968), .Y(n34865) );
  AOI211XL U19051 ( .A0(n34963), .A1(n25127), .B0(n24967), .C0(n24966), .Y(
        n24968) );
  NOR2X1 U19052 ( .A(n24719), .B(n24718), .Y(n24720) );
  NOR2X1 U19053 ( .A(n18379), .B(n18378), .Y(n18380) );
  NAND2XL U19054 ( .A(n25498), .B(n25497), .Y(n34899) );
  AOI211XL U19055 ( .A0(n25766), .A1(n25496), .B0(n25495), .C0(n25494), .Y(
        n25497) );
  NAND2XL U19056 ( .A(n30289), .B(n27736), .Y(n30337) );
  NOR2X1 U19057 ( .A(n27735), .B(n35853), .Y(n30338) );
  NOR2X1 U19058 ( .A(n35853), .B(n27860), .Y(n30332) );
  NOR2X1 U19059 ( .A(n30344), .B(n30343), .Y(n30346) );
  NOR2X1 U19060 ( .A(n35853), .B(n29878), .Y(n29880) );
  NOR2X1 U19061 ( .A(n35853), .B(n19110), .Y(n33056) );
  NAND2XL U19062 ( .A(conv_2[302]), .B(n33057), .Y(n33055) );
  INVXL U19063 ( .A(n33056), .Y(n33058) );
  OAI31XL U19064 ( .A0(n35853), .A1(n31871), .A2(n23856), .B0(n23855), .Y(
        n27412) );
  OAI31XL U19065 ( .A0(n35853), .A1(n28660), .A2(n23708), .B0(n23707), .Y(
        n27051) );
  OAI31XL U19066 ( .A0(n35853), .A1(n22257), .A2(n23350), .B0(n23349), .Y(
        n30414) );
  NAND2XL U19067 ( .A(n35853), .B(n23350), .Y(n23349) );
  ADDFXL U19068 ( .A(conv_2[152]), .B(n24256), .CI(n24255), .CO(n23111), .S(
        n24257) );
  NOR2X1 U19069 ( .A(n35853), .B(n23296), .Y(n24256) );
  OAI31XL U19070 ( .A0(n35853), .A1(n33020), .A2(n23477), .B0(n23476), .Y(
        n30418) );
  OAI31XL U19071 ( .A0(n35853), .A1(n27799), .A2(n23027), .B0(n23026), .Y(
        n31067) );
  NOR2X1 U19072 ( .A(n35853), .B(n35857), .Y(intadd_0_B_0_) );
  NAND2X1 U19073 ( .A(n22896), .B(filter_2_bias[2]), .Y(n34621) );
  NAND4XL U19074 ( .A(n21187), .B(n21186), .C(n21185), .D(n21184), .Y(n35012)
         );
  OAI211XL U19075 ( .A0(n20441), .A1(n25853), .B0(n19495), .C0(n19494), .Y(
        n35024) );
  OAI211XL U19076 ( .A0(n20441), .A1(n34969), .B0(n20440), .C0(n20439), .Y(
        n34976) );
  AOI211XL U19077 ( .A0(n34992), .A1(n21175), .B0(n20438), .C0(n20437), .Y(
        n20439) );
  AOI22XL U19078 ( .A0(N18471), .A1(n26183), .B0(n34963), .B1(n28280), .Y(
        n26186) );
  AOI22XL U19079 ( .A0(n34963), .A1(n35148), .B0(n16671), .B1(n28279), .Y(
        n24838) );
  NOR4XL U19080 ( .A(n28284), .B(n28283), .C(n28282), .D(n28281), .Y(n35007)
         );
  NAND4XL U19081 ( .A(n25723), .B(n25722), .C(n25721), .D(n28275), .Y(n35020)
         );
  NOR2X1 U19082 ( .A(n30536), .B(n27898), .Y(n23954) );
  AOI2BB1XL U19083 ( .A0N(n18997), .A1N(n22269), .B0(n23803), .Y(n35564) );
  INVXL U19084 ( .A(n23219), .Y(n30713) );
  AOI2BB1XL U19085 ( .A0N(n18997), .A1N(n19108), .B0(n23218), .Y(n23219) );
  NOR2X1 U19086 ( .A(n18997), .B(n31871), .Y(n31086) );
  NOR2X1 U19087 ( .A(n30536), .B(n29136), .Y(n22158) );
  NOR2X1 U19088 ( .A(n30742), .B(n30741), .Y(n30744) );
  NAND2X1 U19089 ( .A(n22896), .B(filter_3_bias[2]), .Y(n35566) );
  AOI211XL U19090 ( .A0(conv_1[18]), .A1(n21766), .B0(n21495), .C0(n21494), 
        .Y(n22098) );
  AOI211XL U19091 ( .A0(n16755), .A1(n20214), .B0(n20213), .C0(n20212), .Y(
        n20611) );
  AOI211XL U19092 ( .A0(n28465), .A1(n20214), .B0(n19807), .C0(n19806), .Y(
        n20160) );
  AOI211XL U19093 ( .A0(n26263), .A1(n26385), .B0(n26382), .C0(n25383), .Y(
        n25685) );
  AOI22XL U19094 ( .A0(n28528), .A1(n26537), .B0(n34963), .B1(n25374), .Y(
        n25382) );
  AOI211XL U19095 ( .A0(n28465), .A1(n26389), .B0(n26388), .C0(n26387), .Y(
        n28618) );
  NOR2X1 U19096 ( .A(n24617), .B(n24616), .Y(n34862) );
  ADDFXL U19097 ( .A(conv_1[528]), .B(n32865), .CI(n32864), .CO(n22219), .S(
        n32866) );
  NOR2XL U19098 ( .A(n35498), .B(n33429), .Y(n32865) );
  AOI2BB1XL U19099 ( .A0N(conv_1[527]), .A1N(n30460), .B0(n30461), .Y(n32864)
         );
  AOI2BB1XL U19100 ( .A0N(conv_1[482]), .A1N(n27373), .B0(n27374), .Y(n27224)
         );
  NAND2XL U19101 ( .A(n18851), .B(n26986), .Y(n26951) );
  NOR2X1 U19102 ( .A(n27235), .B(n27234), .Y(n27249) );
  NOR2X1 U19103 ( .A(n29572), .B(n29571), .Y(n29574) );
  ADDFXL U19104 ( .A(conv_1[348]), .B(n24316), .CI(n24315), .CO(n24317), .S(
        n24280) );
  NOR2X1 U19105 ( .A(n24225), .B(n24224), .Y(n24227) );
  NAND2XL U19106 ( .A(n23890), .B(n22295), .Y(n23363) );
  NOR2X1 U19107 ( .A(n23612), .B(n23611), .Y(n23614) );
  NOR2X1 U19108 ( .A(n31370), .B(n31371), .Y(n31369) );
  NOR2X1 U19109 ( .A(n35498), .B(n26509), .Y(n26511) );
  AOI2BB1XL U19110 ( .A0N(conv_1[92]), .A1N(n26684), .B0(n26685), .Y(n26510)
         );
  ADDFXL U19111 ( .A(conv_1[78]), .B(n22867), .CI(n22866), .CO(n22954), .S(
        n22413) );
  NOR2X1 U19112 ( .A(n35498), .B(n33020), .Y(n22867) );
  NAND2X1 U19113 ( .A(n22896), .B(filter_1_bias[3]), .Y(n32867) );
  AOI211XL U19114 ( .A0(n18463), .A1(n25842), .B0(n20977), .C0(n20976), .Y(
        n22051) );
  AOI211XL U19115 ( .A0(n16755), .A1(n25849), .B0(n25848), .C0(n25847), .Y(
        n26118) );
  AOI211XL U19116 ( .A0(n28465), .A1(n25849), .B0(n21825), .C0(n21824), .Y(
        n34873) );
  AOI21XL U19117 ( .A0(N18471), .A1(n25111), .B0(n24963), .Y(n25446) );
  AOI22XL U19118 ( .A0(n16667), .A1(n25104), .B0(n34963), .B1(n25107), .Y(
        n24961) );
  AOI22XL U19119 ( .A0(n28528), .A1(n25104), .B0(n34963), .B1(n25108), .Y(
        n24093) );
  AOI211XL U19120 ( .A0(n26470), .A1(n24707), .B0(n24706), .C0(n24705), .Y(
        n34886) );
  NOR2XL U19121 ( .A(n24702), .B(n35159), .Y(n24706) );
  AOI211XL U19122 ( .A0(n16755), .A1(n24707), .B0(n18364), .C0(n18363), .Y(
        n34942) );
  ADDFXL U19123 ( .A(conv_2[528]), .B(n27685), .CI(n27684), .CO(n27686), .S(
        n24310) );
  NOR2X1 U19124 ( .A(n29644), .B(n29645), .Y(n29643) );
  ADDFXL U19125 ( .A(conv_2[453]), .B(n24338), .CI(n24337), .CO(n27643), .S(
        n23721) );
  NOR2X1 U19126 ( .A(n23992), .B(n23991), .Y(n23994) );
  OAI21XL U19127 ( .A0(n29872), .A1(n29877), .B0(n29873), .Y(n24297) );
  NOR2X1 U19128 ( .A(n28146), .B(n28145), .Y(n23157) );
  NAND2XL U19129 ( .A(n26934), .B(n22961), .Y(n29047) );
  NOR2X1 U19130 ( .A(n35856), .B(n29136), .Y(n29048) );
  NOR2X1 U19131 ( .A(n28652), .B(n28651), .Y(n27083) );
  ADDFXL U19132 ( .A(conv_2[138]), .B(n23038), .CI(n23037), .CO(n22900), .S(
        n23039) );
  NOR2X1 U19133 ( .A(n35856), .B(n34426), .Y(n23038) );
  ADDFXL U19134 ( .A(conv_2[123]), .B(n23334), .CI(n23333), .CO(n23335), .S(
        n23046) );
  NOR2X1 U19135 ( .A(n35856), .B(n28948), .Y(n23334) );
  NOR2X1 U19136 ( .A(n27139), .B(n27140), .Y(n27138) );
  NOR2X1 U19137 ( .A(n26742), .B(n26743), .Y(n26741) );
  NOR2X1 U19138 ( .A(n35856), .B(n35857), .Y(intadd_0_B_1_) );
  NAND2X1 U19139 ( .A(n22896), .B(filter_2_bias[3]), .Y(n34105) );
  NOR4XL U19140 ( .A(n21143), .B(n21142), .C(n21141), .D(n21140), .Y(n35016)
         );
  AOI211XL U19141 ( .A0(n16755), .A1(n20429), .B0(n19469), .C0(n19468), .Y(
        n35028) );
  AOI211XL U19142 ( .A0(n28465), .A1(n20429), .B0(n20428), .C0(n20427), .Y(
        n34980) );
  AOI2BB1XL U19143 ( .A0N(n35126), .A1N(n28479), .B0(n26176), .Y(n34947) );
  AOI22XL U19144 ( .A0(n26263), .A1(n35128), .B0(n34963), .B1(n26170), .Y(
        n26174) );
  AOI21XL U19145 ( .A0(n28465), .A1(n25706), .B0(n18613), .Y(n35019) );
  AOI2BB1XL U19146 ( .A0N(n28274), .A1N(n16701), .B0(n24851), .Y(n24852) );
  OAI21XL U19147 ( .A0(n28274), .A1(n35159), .B0(n28273), .Y(n35008) );
  AOI211XL U19148 ( .A0(n16665), .A1(n35127), .B0(n28272), .C0(n28271), .Y(
        n28273) );
  AOI211XL U19149 ( .A0(n26470), .A1(n25706), .B0(n25705), .C0(n25704), .Y(
        n26704) );
  ADDFXL U19150 ( .A(conv_3[528]), .B(n23735), .CI(n23734), .CO(n23549), .S(
        n23736) );
  NOR2X1 U19151 ( .A(n29426), .B(n33429), .Y(n23735) );
  NOR2X1 U19152 ( .A(n29632), .B(n29631), .Y(n29634) );
  NOR2X1 U19153 ( .A(n29696), .B(n29695), .Y(n29698) );
  NOR2X1 U19154 ( .A(n24203), .B(n24202), .Y(n24205) );
  NOR2X1 U19155 ( .A(n23506), .B(n23505), .Y(n23499) );
  NOR2X1 U19156 ( .A(n29426), .B(n24021), .Y(n29657) );
  NOR2X1 U19157 ( .A(n29657), .B(n29658), .Y(n29656) );
  NOR2X1 U19158 ( .A(n29732), .B(n29733), .Y(n29731) );
  ADDFXL U19159 ( .A(conv_3[168]), .B(n29069), .CI(n29068), .CO(n29071), .S(
        n23750) );
  NOR2X1 U19160 ( .A(n22909), .B(n22908), .Y(n29650) );
  NAND2X1 U19161 ( .A(n22896), .B(filter_3_bias[3]), .Y(n35574) );
  AOI22XL U19162 ( .A0(n26263), .A1(n26412), .B0(n34963), .B1(n25334), .Y(
        n25343) );
  AOI211XL U19163 ( .A0(n26470), .A1(n26416), .B0(n26415), .C0(n26414), .Y(
        n28616) );
  NOR2X1 U19164 ( .A(n24591), .B(n24590), .Y(n24666) );
  INVXL U19165 ( .A(n34860), .Y(n34861) );
  INVXL U19166 ( .A(n34839), .Y(n34835) );
  AOI21XL U19167 ( .A0(n22219), .A1(n22218), .B0(n22220), .Y(n26146) );
  NOR2X1 U19168 ( .A(n27001), .B(n27000), .Y(n27003) );
  AOI2BB1XL U19169 ( .A0N(conv_1[408]), .A1N(n29571), .B0(n29572), .Y(n35483)
         );
  NOR2X1 U19170 ( .A(n35500), .B(n28070), .Y(n35484) );
  NOR2X1 U19171 ( .A(n23760), .B(n23759), .Y(n23762) );
  NOR2X1 U19172 ( .A(n30277), .B(n30276), .Y(n30279) );
  NOR2X1 U19173 ( .A(n30283), .B(n30282), .Y(n30285) );
  ADDFXL U19174 ( .A(conv_1[288]), .B(n24287), .CI(n24286), .CO(n30774), .S(
        n24289) );
  NOR2X1 U19175 ( .A(n35498), .B(n31871), .Y(n24287) );
  AOI2BB1XL U19176 ( .A0N(conv_1[287]), .A1N(n30479), .B0(n30480), .Y(n24286)
         );
  NOR2X1 U19177 ( .A(n35500), .B(n31871), .Y(n30773) );
  NOR2X1 U19178 ( .A(n30773), .B(n30774), .Y(n30772) );
  ADDFXL U19179 ( .A(conv_1[273]), .B(n22387), .CI(n22386), .CO(n30767), .S(
        n22388) );
  NOR2X1 U19180 ( .A(n35498), .B(n33994), .Y(n22387) );
  AOI2BB1XL U19181 ( .A0N(conv_1[272]), .A1N(n30473), .B0(n30474), .Y(n22386)
         );
  NOR2X1 U19182 ( .A(n35500), .B(n33994), .Y(n30766) );
  NOR2X1 U19183 ( .A(n30766), .B(n30767), .Y(n30765) );
  NOR2X1 U19184 ( .A(n24692), .B(n24691), .Y(n33215) );
  AND2XL U19185 ( .A(n24692), .B(n24691), .Y(n33219) );
  NOR2X1 U19186 ( .A(n24439), .B(n24440), .Y(n24438) );
  NOR2X1 U19187 ( .A(n24169), .B(n24168), .Y(n24171) );
  NOR2X1 U19188 ( .A(n23976), .B(n23975), .Y(n23978) );
  NOR2X1 U19189 ( .A(n24496), .B(n24497), .Y(n24495) );
  NOR2X1 U19190 ( .A(n24008), .B(n24009), .Y(n24007) );
  NOR2X1 U19191 ( .A(n30754), .B(n30753), .Y(n30756) );
  NOR2X1 U19192 ( .A(n26922), .B(n26921), .Y(n26924) );
  NOR2X1 U19193 ( .A(n27405), .B(n27406), .Y(n27404) );
  NOR2X1 U19194 ( .A(n27037), .B(n27036), .Y(n27039) );
  NAND2X1 U19195 ( .A(n22896), .B(filter_1_bias[4]), .Y(n35489) );
  NOR4XL U19196 ( .A(n20794), .B(n20793), .C(n20792), .D(n20791), .Y(n22053)
         );
  AOI22XL U19197 ( .A0(n34963), .A1(n25134), .B0(n26172), .B1(n25501), .Y(
        n24980) );
  AOI211XL U19198 ( .A0(n34963), .A1(n25135), .B0(n24058), .C0(n24057), .Y(
        n24059) );
  AOI22XL U19199 ( .A0(n34963), .A1(n25132), .B0(n28324), .B1(n25135), .Y(
        n24725) );
  INVXL U19200 ( .A(n34940), .Y(n34943) );
  NOR2X1 U19201 ( .A(n28853), .B(n28852), .Y(n28855) );
  NOR2X1 U19202 ( .A(n28990), .B(n28989), .Y(n28992) );
  NOR2X1 U19203 ( .A(n28984), .B(n28983), .Y(n28986) );
  NOR2X1 U19204 ( .A(n28075), .B(n28074), .Y(n28858) );
  AOI2BB1XL U19205 ( .A0N(conv_2[393]), .A1N(n29565), .B0(n29566), .Y(n29055)
         );
  NOR2X1 U19206 ( .A(n35858), .B(n32016), .Y(n29056) );
  NOR2X1 U19207 ( .A(n24192), .B(n24193), .Y(n24191) );
  NOR2X1 U19208 ( .A(n28865), .B(n28864), .Y(n28867) );
  NOR2X1 U19209 ( .A(n28871), .B(n28870), .Y(n28873) );
  NOR2X1 U19210 ( .A(n29062), .B(n29063), .Y(n29061) );
  NOR2X1 U19211 ( .A(n35856), .B(n28721), .Y(n32984) );
  NOR2X1 U19212 ( .A(n35858), .B(n28721), .Y(n29408) );
  NOR2X1 U19213 ( .A(n29408), .B(n29409), .Y(n29407) );
  NOR2X1 U19214 ( .A(n28148), .B(n28147), .Y(n28977) );
  NOR2X1 U19215 ( .A(n29050), .B(n29049), .Y(n29138) );
  NOR2X1 U19216 ( .A(n29023), .B(n29022), .Y(n29025) );
  NOR2X1 U19217 ( .A(n23370), .B(n23369), .Y(n23372) );
  NOR2X1 U19218 ( .A(n27970), .B(n27971), .Y(n22903) );
  NOR2X1 U19219 ( .A(n24352), .B(n24353), .Y(n23338) );
  NOR2X1 U19220 ( .A(n24015), .B(n24016), .Y(n24014) );
  NOR2X1 U19221 ( .A(n28740), .B(n28741), .Y(n23482) );
  NOR2X1 U19222 ( .A(n29739), .B(n29740), .Y(n29738) );
  NAND2X1 U19223 ( .A(n22896), .B(filter_2_bias[4]), .Y(n34408) );
  NOR4BXL U19224 ( .AN(n21210), .B(n21209), .C(n21208), .D(n21207), .Y(n22107)
         );
  INVXL U19225 ( .A(n34978), .Y(n34979) );
  AOI211XL U19226 ( .A0(n16667), .A1(n35102), .B0(n26212), .C0(n26211), .Y(
        n27067) );
  AOI22XL U19227 ( .A0(n26263), .A1(n35101), .B0(n34963), .B1(n26208), .Y(
        n26209) );
  INVXL U19228 ( .A(n35250), .Y(n35252) );
  NOR2X1 U19229 ( .A(n24364), .B(n24365), .Y(n23552) );
  NOR2X1 U19230 ( .A(n23772), .B(n23773), .Y(n23519) );
  ADDFXL U19231 ( .A(conv_3[453]), .B(n23049), .CI(n23048), .CO(n24261), .S(
        n23050) );
  NOR2X1 U19232 ( .A(n27644), .B(n29426), .Y(n23049) );
  NOR2X1 U19233 ( .A(n24260), .B(n24261), .Y(n24259) );
  NOR2X1 U19234 ( .A(n31925), .B(n31926), .Y(n23962) );
  NOR2X1 U19235 ( .A(n26814), .B(n26815), .Y(n26813) );
  NOR2X1 U19236 ( .A(n31625), .B(n31626), .Y(n23511) );
  NOR2X1 U19237 ( .A(n31392), .B(n31391), .Y(n26718) );
  OAI2BB1XL U19238 ( .A0N(conv_3[318]), .A1N(n23811), .B0(n23810), .Y(n28755)
         );
  NOR2X1 U19239 ( .A(n31691), .B(n28721), .Y(n28723) );
  NOR2X1 U19240 ( .A(n22146), .B(n22145), .Y(n24474) );
  NOR2X1 U19241 ( .A(n26315), .B(n26316), .Y(n22135) );
  NOR2BXL U19242 ( .AN(n29072), .B(conv_3[169]), .Y(n31560) );
  NOR2X1 U19243 ( .A(n28949), .B(n28950), .Y(n23692) );
  NOR2X1 U19244 ( .A(n22911), .B(n22910), .Y(n31768) );
  NOR2X1 U19245 ( .A(n31803), .B(n31804), .Y(n22923) );
  NOR2X1 U19246 ( .A(n24469), .B(n24468), .Y(n29663) );
  NOR2X1 U19247 ( .A(n30196), .B(n30197), .Y(n29434) );
  NAND2X1 U19248 ( .A(n22896), .B(filter_3_bias[4]), .Y(n34097) );
  NOR2XL U19249 ( .A(n29216), .B(n26965), .Y(n26964) );
  ADDFXL U19250 ( .A(conv_1[536]), .B(n29216), .CI(n26960), .CO(n26965), .S(
        n22223) );
  AOI2BB1XL U19251 ( .A0N(conv_1[535]), .A1N(n29189), .B0(n29190), .Y(n26960)
         );
  NOR2X1 U19252 ( .A(n29190), .B(n29189), .Y(n29192) );
  AOI2BB1XL U19253 ( .A0N(conv_1[533]), .A1N(n29234), .B0(n29236), .Y(n29214)
         );
  OAI32XL U19254 ( .A0(n29236), .A1(conv_1[530]), .A2(n23696), .B0(n29216), 
        .B1(n22221), .Y(n29242) );
  NAND2XL U19255 ( .A(n29242), .B(conv_1[531]), .Y(n29241) );
  NOR4XL U19256 ( .A(n21477), .B(n21476), .C(n21475), .D(n21474), .Y(n21793)
         );
  OAI21XL U19257 ( .A0(n35229), .A1(n21791), .B0(n35227), .Y(n34815) );
  AOI222XL U19258 ( .A0(n21790), .A1(n21789), .B0(n21790), .B1(n21788), .C0(
        n21789), .C1(n21787), .Y(n21791) );
  AOI211XL U19259 ( .A0(n16755), .A1(n20193), .B0(n20192), .C0(n20191), .Y(
        n20351) );
  OAI211XL U19260 ( .A0(n36246), .A1(n25297), .B0(n16659), .C0(n20185), .Y(
        n20186) );
  AOI21XL U19261 ( .A0(n35227), .A1(n20349), .B0(n28595), .Y(n34844) );
  AOI222XL U19262 ( .A0(n20348), .A1(n20347), .B0(n20348), .B1(n20346), .C0(
        n20347), .C1(n20345), .Y(n20349) );
  AOI22XL U19263 ( .A0(n34963), .A1(n21467), .B0(n35234), .B1(n21458), .Y(
        n19760) );
  OAI21XL U19264 ( .A0(n35229), .A1(n20099), .B0(n35227), .Y(n34800) );
  AOI21XL U19265 ( .A0(n35227), .A1(n28596), .B0(n28595), .Y(n34821) );
  AOI222XL U19266 ( .A0(n28594), .A1(n28593), .B0(n28594), .B1(n28592), .C0(
        n28593), .C1(n28591), .Y(n28596) );
  AOI211XL U19267 ( .A0(n26470), .A1(n26381), .B0(n26380), .C0(n26379), .Y(
        n26493) );
  OAI21XL U19268 ( .A0(n35229), .A1(n26491), .B0(n35227), .Y(n34806) );
  AOI222XL U19269 ( .A0(n26490), .A1(n26489), .B0(n26490), .B1(n26488), .C0(
        n26489), .C1(n26487), .Y(n26491) );
  NOR4XL U19270 ( .A(n26536), .B(n26535), .C(n26534), .D(n26533), .Y(n26666)
         );
  OAI21XL U19271 ( .A0(n35229), .A1(n26664), .B0(n35227), .Y(n34810) );
  AOI222XL U19272 ( .A0(n26663), .A1(n26662), .B0(n26663), .B1(n26661), .C0(
        n26662), .C1(n26660), .Y(n26664) );
  INVX2 U19273 ( .A(n18535), .Y(n26621) );
  AOI2BB2XL U19274 ( .B0(n30267), .B1(n25261), .A0N(n25262), .A1N(n25260), .Y(
        n30262) );
  NAND2XL U19275 ( .A(n30262), .B(conv_1[519]), .Y(n30266) );
  NAND2XL U19276 ( .A(n25259), .B(n25261), .Y(n27257) );
  NAND2XL U19277 ( .A(n27131), .B(n27114), .Y(n27133) );
  NOR2X1 U19278 ( .A(n27124), .B(n27118), .Y(n27126) );
  AOI21XL U19279 ( .A0(n26339), .A1(n26334), .B0(n23427), .Y(n23653) );
  NOR2X1 U19280 ( .A(n27131), .B(n26335), .Y(n23427) );
  AOI2BB1XL U19281 ( .A0N(conv_1[488]), .A1N(n35539), .B0(n35534), .Y(n29982)
         );
  AOI2BB1XL U19282 ( .A0N(conv_1[486]), .A1N(n35526), .B0(n35534), .Y(n35532)
         );
  AOI2BB1XL U19283 ( .A0N(conv_1[485]), .A1N(n29971), .B0(n35534), .Y(n35526)
         );
  NOR2X1 U19284 ( .A(n27603), .B(n27604), .Y(n27173) );
  AOI2BB1XL U19285 ( .A0N(conv_1[471]), .A1N(n27178), .B0(n29823), .Y(n27602)
         );
  INVXL U19286 ( .A(n32887), .Y(n29823) );
  NOR2X1 U19287 ( .A(n33161), .B(n29823), .Y(n27178) );
  NOR2X1 U19288 ( .A(n33166), .B(n20008), .Y(n27179) );
  AND2XL U19289 ( .A(n32887), .B(n18855), .Y(n33162) );
  NOR2X1 U19290 ( .A(n27860), .B(n18847), .Y(n33507) );
  INVXL U19291 ( .A(n27860), .Y(n33509) );
  OAI2BB1XL U19292 ( .A0N(conv_1[461]), .A1N(n30024), .B0(n30051), .Y(n28729)
         );
  NOR2X1 U19293 ( .A(conv_1[461]), .B(n30025), .Y(n28731) );
  OAI2BB1XL U19294 ( .A0N(conv_1[460]), .A1N(n30043), .B0(n30051), .Y(n30024)
         );
  OR2XL U19295 ( .A(n30051), .B(n27239), .Y(n30042) );
  AOI2BB1XL U19296 ( .A0N(conv_1[456]), .A1N(n30018), .B0(n30051), .Y(n30049)
         );
  AOI2BB1XL U19297 ( .A0N(conv_1[455]), .A1N(n27244), .B0(n30051), .Y(n30018)
         );
  NOR2X1 U19298 ( .A(n27243), .B(n27248), .Y(n30019) );
  INVXL U19299 ( .A(n30051), .Y(n30044) );
  NOR2X1 U19300 ( .A(n33423), .B(n27644), .Y(n27422) );
  NAND2XL U19301 ( .A(n27422), .B(conv_1[450]), .Y(n27421) );
  NOR2BXL U19302 ( .AN(n35521), .B(conv_1[446]), .Y(n35523) );
  OAI2BB1XL U19303 ( .A0N(conv_1[445]), .A1N(n35514), .B0(n27149), .Y(n35522)
         );
  AOI2BB1XL U19304 ( .A0N(conv_1[444]), .A1N(n27161), .B0(n27149), .Y(n35513)
         );
  NOR2X1 U19305 ( .A(n35515), .B(n27161), .Y(n27160) );
  ADDFXL U19306 ( .A(conv_1[443]), .B(n35515), .CI(n27145), .CO(n27161), .S(
        n23644) );
  AOI21XL U19307 ( .A0(n25231), .A1(n25236), .B0(n25232), .Y(n27145) );
  NOR2X1 U19308 ( .A(n29223), .B(n29222), .Y(n35508) );
  NOR2X1 U19309 ( .A(conv_1[429]), .B(n33392), .Y(n33393) );
  NOR2X1 U19310 ( .A(n27585), .B(n27584), .Y(n33394) );
  NOR2X1 U19311 ( .A(n27582), .B(n29328), .Y(n33392) );
  NOR2X1 U19312 ( .A(intadd_1_B_2_), .B(n33394), .Y(n33391) );
  NOR2X1 U19313 ( .A(n27594), .B(n34775), .Y(n33385) );
  NOR2X1 U19314 ( .A(n35493), .B(n33387), .Y(n33384) );
  AOI2BB1XL U19315 ( .A0N(conv_1[412]), .A1N(n35491), .B0(n34775), .Y(n27595)
         );
  NOR2X1 U19316 ( .A(conv_1[413]), .B(n27595), .Y(n27594) );
  AOI2BB1XL U19317 ( .A0N(conv_1[411]), .A1N(n29286), .B0(n34775), .Y(n35491)
         );
  NOR2X1 U19318 ( .A(n29287), .B(n29291), .Y(n35492) );
  NOR2X1 U19319 ( .A(n29357), .B(n29356), .Y(n31279) );
  AOI2BB1XL U19320 ( .A0N(conv_1[396]), .A1N(n29268), .B0(n35471), .Y(n27639)
         );
  AOI2BB1XL U19321 ( .A0N(conv_1[395]), .A1N(n29275), .B0(n35471), .Y(n29268)
         );
  NOR2X1 U19322 ( .A(n29274), .B(n29279), .Y(n29269) );
  AOI21XL U19323 ( .A0(n34340), .A1(n34335), .B0(n34336), .Y(n22975) );
  AOI2BB1XL U19324 ( .A0N(conv_1[382]), .A1N(n23128), .B0(n33088), .Y(n35461)
         );
  NOR2X1 U19325 ( .A(n23129), .B(n23133), .Y(n35462) );
  AOI2BB1XL U19326 ( .A0N(conv_1[381]), .A1N(n23134), .B0(n33088), .Y(n23128)
         );
  INVXL U19327 ( .A(n35463), .Y(n33088) );
  NOR2BXL U19328 ( .AN(conv_1[380]), .B(n33181), .Y(n23135) );
  AND2XL U19329 ( .A(n35463), .B(n19153), .Y(n33177) );
  NOR2X1 U19330 ( .A(n27578), .B(n27577), .Y(n35454) );
  NAND2XL U19331 ( .A(conv_1[360]), .B(n30058), .Y(n30057) );
  INVXL U19332 ( .A(n35441), .Y(n28847) );
  NOR2BXL U19333 ( .AN(n35448), .B(conv_1[356]), .Y(n35450) );
  OAI2BB1XL U19334 ( .A0N(conv_1[355]), .A1N(n28815), .B0(n28847), .Y(n35449)
         );
  AOI2BB1XL U19335 ( .A0N(conv_1[354]), .A1N(n35442), .B0(n28847), .Y(n28816)
         );
  NOR2X1 U19336 ( .A(n35440), .B(n35444), .Y(n28815) );
  ADDFXL U19337 ( .A(conv_1[353]), .B(n35441), .CI(n28804), .CO(n35442), .S(
        n24320) );
  AOI2BB1XL U19338 ( .A0N(conv_1[352]), .A1N(n28809), .B0(n28810), .Y(n28804)
         );
  AOI2BB1XL U19339 ( .A0N(conv_1[350]), .A1N(n26363), .B0(n28847), .Y(n33643)
         );
  NOR2X1 U19340 ( .A(n35441), .B(n33645), .Y(n33642) );
  NOR2X1 U19341 ( .A(n23015), .B(n23011), .Y(n23005) );
  AOI2BB1XL U19342 ( .A0N(conv_1[338]), .A1N(n35432), .B0(n28821), .Y(n23010)
         );
  NOR2X1 U19343 ( .A(n23000), .B(n22999), .Y(n35433) );
  ADDFXL U19344 ( .A(conv_1[334]), .B(n24241), .CI(n24240), .CO(n22994), .S(
        n24243) );
  AOI2BB1XL U19345 ( .A0N(conv_1[333]), .A1N(n23140), .B0(n23141), .Y(n24240)
         );
  NOR2X1 U19346 ( .A(n35434), .B(n22994), .Y(n22988) );
  NOR2X1 U19347 ( .A(n34522), .B(n34521), .Y(n34523) );
  ADDFXL U19348 ( .A(conv_1[311]), .B(n28644), .CI(n24158), .CO(n24175), .S(
        n22320) );
  AOI21XL U19349 ( .A0(n25282), .A1(n25287), .B0(n25283), .Y(n24158) );
  OAI2BB1XL U19350 ( .A0N(n28643), .A1N(conv_1[308]), .B0(n24159), .Y(n24163)
         );
  NAND2XL U19351 ( .A(n22549), .B(n28646), .Y(n28649) );
  NAND2XL U19352 ( .A(n28644), .B(n22317), .Y(n28646) );
  AOI2BB1XL U19353 ( .A0N(n24153), .A1N(conv_1[306]), .B0(n24159), .Y(n19218)
         );
  NOR2X1 U19354 ( .A(n28644), .B(n24153), .Y(n24152) );
  NOR2X1 U19355 ( .A(n22826), .B(n23169), .Y(n23176) );
  NOR2BXL U19356 ( .AN(n35421), .B(conv_1[278]), .Y(n35423) );
  OAI2BB1XL U19357 ( .A0N(n29345), .A1N(conv_1[277]), .B0(n29339), .Y(n35422)
         );
  AOI2BB1XL U19358 ( .A0N(conv_1[275]), .A1N(n29370), .B0(n29339), .Y(n29316)
         );
  NOR2X1 U19359 ( .A(n33663), .B(n35411), .Y(n23836) );
  ADDFXL U19360 ( .A(conv_1[247]), .B(n33663), .CI(n23659), .CO(n23835), .S(
        n22312) );
  AOI21XL U19361 ( .A0(n34333), .A1(n34328), .B0(n34329), .Y(n23659) );
  NOR2X1 U19362 ( .A(n35414), .B(n22311), .Y(n23841) );
  AOI2BB1XL U19363 ( .A0N(n35404), .A1N(n31128), .B0(n31127), .Y(n26674) );
  ADDFXL U19364 ( .A(conv_1[233]), .B(n35404), .CI(n26672), .CO(n35405), .S(
        n22300) );
  NOR2BXL U19365 ( .AN(n35399), .B(n35400), .Y(n26672) );
  NOR2BXL U19366 ( .AN(n35398), .B(conv_1[232]), .Y(n35400) );
  OAI2BB1XL U19367 ( .A0N(n29263), .A1N(conv_1[231]), .B0(n34276), .Y(n35399)
         );
  NOR2X1 U19368 ( .A(n33182), .B(n34276), .Y(n29262) );
  NOR2X1 U19369 ( .A(n33187), .B(n22571), .Y(n29263) );
  AND2XL U19370 ( .A(n35404), .B(n22299), .Y(n33183) );
  NOR2X1 U19371 ( .A(n29136), .B(n22291), .Y(n33873) );
  AOI2BB1XL U19372 ( .A0N(conv_1[216]), .A1N(n23303), .B0(n28602), .Y(n35390)
         );
  NOR2X1 U19373 ( .A(n23308), .B(n23304), .Y(n35391) );
  AOI2BB1XL U19374 ( .A0N(conv_1[215]), .A1N(n23341), .B0(n28602), .Y(n23303)
         );
  NOR2X1 U19375 ( .A(n28660), .B(n23286), .Y(n33869) );
  AOI2BB1XL U19376 ( .A0N(conv_1[204]), .A1N(n31113), .B0(n34060), .Y(n35377)
         );
  NOR2X1 U19377 ( .A(n31112), .B(n31111), .Y(n35378) );
  AOI2BB1XL U19378 ( .A0N(conv_1[203]), .A1N(n35371), .B0(n34060), .Y(n31113)
         );
  AOI2BB1XL U19379 ( .A0N(conv_1[202]), .A1N(n23451), .B0(n34060), .Y(n35371)
         );
  NOR2X1 U19380 ( .A(n23450), .B(n23449), .Y(n35372) );
  NOR2X1 U19381 ( .A(n23681), .B(n34060), .Y(n23451) );
  NOR2X1 U19382 ( .A(n33423), .B(n27848), .Y(n24217) );
  AOI2BB1XL U19383 ( .A0N(conv_1[186]), .A1N(n35351), .B0(n32988), .Y(n23599)
         );
  NOR2X1 U19384 ( .A(n33188), .B(n32988), .Y(n35351) );
  NOR2X1 U19385 ( .A(n33193), .B(n23592), .Y(n35352) );
  AND2XL U19386 ( .A(n35365), .B(n23593), .Y(n33189) );
  NOR2X1 U19387 ( .A(n33423), .B(n34703), .Y(n24138) );
  NAND2XL U19388 ( .A(n24138), .B(conv_1[180]), .Y(n24137) );
  ADDFXL U19389 ( .A(conv_1[176]), .B(n23923), .CI(n23916), .CO(n26667), .S(
        n22303) );
  ADDFXL U19390 ( .A(conv_1[175]), .B(n23923), .CI(n22302), .CO(n23916), .S(
        n22281) );
  AOI2BB1XL U19391 ( .A0N(conv_1[174]), .A1N(n23935), .B0(n23936), .Y(n22302)
         );
  AND2XL U19392 ( .A(n27543), .B(n27542), .Y(n27540) );
  NOR2BXL U19393 ( .AN(n35347), .B(n35348), .Y(n22280) );
  OAI2BB1XL U19394 ( .A0N(n26671), .A1N(n29676), .B0(n24673), .Y(n23915) );
  NOR2X1 U19395 ( .A(conv_1[170]), .B(n35344), .Y(n35348) );
  NOR2X1 U19396 ( .A(n22257), .B(n22258), .Y(n33497) );
  NAND2XL U19397 ( .A(n34044), .B(n23299), .Y(n23376) );
  NOR2X1 U19398 ( .A(n23398), .B(n23393), .Y(n23388) );
  NOR2X1 U19399 ( .A(n23406), .B(n23405), .Y(n23408) );
  NOR2X1 U19400 ( .A(n33423), .B(n23296), .Y(n26691) );
  NOR2X1 U19401 ( .A(conv_1[147]), .B(n32784), .Y(n32781) );
  AOI2BB1XL U19402 ( .A0N(conv_1[143]), .A1N(n26765), .B0(n26766), .Y(n22277)
         );
  NOR2X1 U19403 ( .A(n26766), .B(n26765), .Y(n26768) );
  AOI2BB1XL U19404 ( .A0N(conv_1[141]), .A1N(n26760), .B0(n32780), .Y(n35337)
         );
  NOR2X1 U19405 ( .A(n26759), .B(n26764), .Y(n35338) );
  NOR2X1 U19406 ( .A(n34426), .B(n33501), .Y(n33502) );
  AND2XL U19407 ( .A(n27548), .B(n27547), .Y(n30451) );
  AOI2BB1XL U19408 ( .A0N(conv_1[125]), .A1N(n29304), .B0(n29305), .Y(n23656)
         );
  NOR2X1 U19409 ( .A(n29305), .B(n29304), .Y(n29307) );
  AOI2BB1XL U19410 ( .A0N(conv_1[99]), .A1N(n26797), .B0(n31334), .Y(n26802)
         );
  NOR2X1 U19411 ( .A(n26796), .B(n26795), .Y(n26803) );
  AOI2BB1XL U19412 ( .A0N(conv_1[97]), .A1N(n26807), .B0(n31334), .Y(n26783)
         );
  NOR2X1 U19413 ( .A(n26812), .B(n26808), .Y(n26784) );
  NOR2X1 U19414 ( .A(n34053), .B(n26724), .Y(n26723) );
  ADDFXL U19415 ( .A(conv_1[84]), .B(n34053), .CI(n24926), .CO(n26724), .S(
        n24343) );
  AOI21XL U19416 ( .A0(n24919), .A1(n24924), .B0(n24920), .Y(n24926) );
  NOR2X1 U19417 ( .A(n33020), .B(n22408), .Y(n33494) );
  NOR2X1 U19418 ( .A(n27089), .B(n27088), .Y(n27091) );
  AOI2BB1XL U19419 ( .A0N(conv_1[65]), .A1N(n27107), .B0(n35324), .Y(n27100)
         );
  NOR2X1 U19420 ( .A(n27106), .B(n27111), .Y(n27101) );
  NOR2XL U19421 ( .A(n31418), .B(n22416), .Y(n33488) );
  AOI2BB1XL U19422 ( .A0N(conv_1[54]), .A1N(n35307), .B0(n35309), .Y(n35314)
         );
  NOR2X1 U19423 ( .A(n35311), .B(n35308), .Y(n35315) );
  INVXL U19424 ( .A(n35309), .Y(n35316) );
  AOI2BB1XL U19425 ( .A0N(conv_1[51]), .A1N(n26134), .B0(n35309), .Y(n26820)
         );
  AOI21XL U19426 ( .A0(n35309), .A1(n27322), .B0(n26134), .Y(n27313) );
  MXI2XL U19427 ( .A(n35309), .B(n35316), .S0(n26133), .Y(n27323) );
  NOR3XL U19428 ( .A(n33514), .B(n33423), .C(n27799), .Y(n33512) );
  AOI2BB1XL U19429 ( .A0N(conv_1[38]), .A1N(n27300), .B0(n35289), .Y(n27306)
         );
  NOR2X1 U19430 ( .A(n35288), .B(n35291), .Y(n27301) );
  AOI2BB1XL U19431 ( .A0N(conv_1[35]), .A1N(n27294), .B0(n35289), .Y(n35281)
         );
  NOR2X1 U19432 ( .A(n27295), .B(n27299), .Y(n35282) );
  ADDFXL U19433 ( .A(conv_1[42]), .B(n35296), .CI(n33123), .CO(n33251), .S(
        n25081) );
  NOR2BXL U19434 ( .AN(n35303), .B(n35304), .Y(n33123) );
  NOR2X1 U19435 ( .A(n27343), .B(n27339), .Y(n27351) );
  AOI2BB1XL U19436 ( .A0N(conv_1[21]), .A1N(n27344), .B0(n30588), .Y(n27338)
         );
  AOI2BB1XL U19437 ( .A0N(conv_1[20]), .A1N(n27332), .B0(n30588), .Y(n27344)
         );
  NOR2X1 U19438 ( .A(n27334), .B(n27333), .Y(n27345) );
  NOR2X1 U19439 ( .A(n27278), .B(n27279), .Y(n27277) );
  OAI2BB1XL U19440 ( .A0N(n27285), .A1N(conv_1[7]), .B0(n22380), .Y(n22383) );
  NOR2X1 U19441 ( .A(intadd_2_n1), .B(conv_1[5]), .Y(n27076) );
  NAND2X1 U19442 ( .A(n22896), .B(filter_1_bias[0]), .Y(n34773) );
  NOR2X1 U19443 ( .A(conv_2[536]), .B(n29101), .Y(n28254) );
  NOR2X1 U19444 ( .A(n28254), .B(n29100), .Y(n28252) );
  AOI2BB1XL U19445 ( .A0N(conv_2[532]), .A1N(n29087), .B0(n29095), .Y(n33626)
         );
  NOR2X1 U19446 ( .A(n33629), .B(n33628), .Y(n33625) );
  NOR2X1 U19447 ( .A(conv_2[533]), .B(n33626), .Y(n33627) );
  NOR2X1 U19448 ( .A(n29092), .B(n29088), .Y(n33628) );
  AOI2BB1XL U19449 ( .A0N(conv_2[531]), .A1N(n29625), .B0(n29095), .Y(n29087)
         );
  INVXL U19450 ( .A(n33629), .Y(n29095) );
  OR2X1 U19451 ( .A(n16760), .B(n21810), .Y(n21729) );
  NAND2XL U19452 ( .A(n23055), .B(n16706), .Y(n21730) );
  OAI21XL U19453 ( .A0(n35229), .A1(n21089), .B0(n35227), .Y(n34890) );
  AOI222XL U19454 ( .A0(n21088), .A1(n21087), .B0(n21088), .B1(n21086), .C0(
        n21087), .C1(n21085), .Y(n21089) );
  BUFX2 U19455 ( .A(n16708), .Y(n35159) );
  NAND2X1 U19456 ( .A(n19221), .B(n28467), .Y(n16708) );
  NAND2X1 U19457 ( .A(n36244), .B(n16755), .Y(n26409) );
  NOR2X1 U19458 ( .A(n34904), .B(n20742), .Y(n21801) );
  AOI22XL U19459 ( .A0(n34963), .A1(n34914), .B0(n35234), .B1(n34912), .Y(
        n21806) );
  OAI21XL U19460 ( .A0(n35229), .A1(n22047), .B0(n35227), .Y(n34871) );
  AOI21XL U19461 ( .A0(N18471), .A1(n25103), .B0(n24955), .Y(n25061) );
  AOI22XL U19462 ( .A0(n34992), .A1(n34930), .B0(n34963), .B1(n25100), .Y(
        n24952) );
  OAI21XL U19463 ( .A0(n35229), .A1(n25059), .B0(n35227), .Y(n34866) );
  AOI222XL U19464 ( .A0(n25058), .A1(n25057), .B0(n25058), .B1(n25056), .C0(
        n25057), .C1(n25055), .Y(n25059) );
  AOI21XL U19465 ( .A0(n35227), .A1(n25228), .B0(n28595), .Y(n34896) );
  AOI222XL U19466 ( .A0(n25227), .A1(n25226), .B0(n25227), .B1(n25225), .C0(
        n25226), .C1(n25224), .Y(n25228) );
  AOI211XL U19467 ( .A0(n26470), .A1(n34927), .B0(n24051), .C0(n24050), .Y(
        n24136) );
  OAI21XL U19468 ( .A0(n35229), .A1(n24134), .B0(n35227), .Y(n34880) );
  AOI222XL U19469 ( .A0(n24133), .A1(n24132), .B0(n24133), .B1(n24131), .C0(
        n24132), .C1(n24130), .Y(n24134) );
  AOI211XL U19470 ( .A0(n34927), .A1(n34827), .B0(n24701), .C0(n24700), .Y(
        n24807) );
  AOI22XL U19471 ( .A0(n34963), .A1(n25098), .B0(n28366), .B1(n34930), .Y(
        n24699) );
  OAI21XL U19472 ( .A0(n35229), .A1(n24805), .B0(n35227), .Y(n34884) );
  AOI222XL U19473 ( .A0(n24804), .A1(n24803), .B0(n24804), .B1(n24802), .C0(
        n24803), .C1(n24801), .Y(n24805) );
  OAI211XL U19474 ( .A0(n26575), .A1(n24783), .B0(n24782), .C0(n24781), .Y(
        n24803) );
  NOR2X1 U19475 ( .A(n25466), .B(n25465), .Y(n25674) );
  OAI21XL U19476 ( .A0(n35229), .A1(n25672), .B0(n35227), .Y(n34901) );
  AOI222XL U19477 ( .A0(n25671), .A1(n25670), .B0(n25671), .B1(n25669), .C0(
        n25670), .C1(n25668), .Y(n25672) );
  NOR2X1 U19478 ( .A(n33578), .B(n28706), .Y(n27787) );
  NOR2X1 U19479 ( .A(n33580), .B(n33579), .Y(n33576) );
  NOR2X1 U19480 ( .A(n27775), .B(n27780), .Y(n33579) );
  NAND2XL U19481 ( .A(conv_2[510]), .B(n23253), .Y(n23565) );
  NOR2X1 U19482 ( .A(conv_2[507]), .B(n33172), .Y(n33705) );
  AND2XL U19483 ( .A(n33168), .B(n33167), .Y(n33169) );
  AOI2BB1XL U19484 ( .A0N(conv_2[504]), .A1N(n36079), .B0(n36081), .Y(n36086)
         );
  AOI2BB1XL U19485 ( .A0N(conv_2[503]), .A1N(n36073), .B0(n36081), .Y(n36079)
         );
  NAND2XL U19486 ( .A(n33424), .B(n28739), .Y(n36081) );
  AOI21XL U19487 ( .A0(conv_2[501]), .A1(n27910), .B0(n36088), .Y(n30911) );
  NAND2BXL U19488 ( .AN(conv_2[501]), .B(n18938), .Y(n30909) );
  OR2XL U19489 ( .A(n36081), .B(n18936), .Y(n18938) );
  NOR2X1 U19490 ( .A(n31017), .B(n31016), .Y(n31019) );
  NAND2XL U19491 ( .A(n36088), .B(n33705), .Y(n34011) );
  ADDFXL U19492 ( .A(conv_2[491]), .B(n34132), .CI(n33667), .CO(n34133), .S(
        n29579) );
  AOI2BB1XL U19493 ( .A0N(conv_2[490]), .A1N(n29578), .B0(n29577), .Y(n33667)
         );
  NOR2X1 U19494 ( .A(n34132), .B(n27753), .Y(n27752) );
  NOR2X1 U19495 ( .A(n27759), .B(n27758), .Y(n27761) );
  AOI2BB1XL U19496 ( .A0N(conv_2[485]), .A1N(n27745), .B0(n34130), .Y(n33600)
         );
  NOR2X1 U19497 ( .A(n34132), .B(n33602), .Y(n33599) );
  NOR2X1 U19498 ( .A(conv_2[486]), .B(n33600), .Y(n33601) );
  NOR2X1 U19499 ( .A(n27747), .B(n27746), .Y(n33602) );
  NOR2X1 U19500 ( .A(n27735), .B(n33989), .Y(n23799) );
  NAND2XL U19501 ( .A(n23799), .B(conv_2[480]), .Y(n27734) );
  NAND3BXL U19502 ( .AN(n34133), .B(n34132), .C(n34131), .Y(n34663) );
  NOR2X1 U19503 ( .A(n27891), .B(n27896), .Y(n27944) );
  OR2XL U19504 ( .A(n27943), .B(n27874), .Y(n27885) );
  NOR2X1 U19505 ( .A(n33989), .B(n27860), .Y(n22886) );
  NOR2X1 U19506 ( .A(conv_2[461]), .B(n27660), .Y(n27680) );
  NOR2X1 U19507 ( .A(n27680), .B(n27661), .Y(n27678) );
  AOI2BB1XL U19508 ( .A0N(conv_2[459]), .A1N(n27653), .B0(n27677), .Y(n33608)
         );
  NOR2X1 U19509 ( .A(n33611), .B(n33610), .Y(n33607) );
  OAI21XL U19510 ( .A0(conv_2[457]), .A1(n27666), .B0(n33611), .Y(n27671) );
  NOR2X1 U19511 ( .A(n33611), .B(n30876), .Y(n27645) );
  NOR2X1 U19512 ( .A(n27644), .B(n23716), .Y(n34442) );
  AOI2BB1XL U19513 ( .A0N(conv_2[444]), .A1N(n28790), .B0(n28937), .Y(n27922)
         );
  AOI2BB1XL U19514 ( .A0N(conv_2[443]), .A1N(n36065), .B0(n28937), .Y(n28790)
         );
  AOI2BB1XL U19515 ( .A0N(conv_2[441]), .A1N(n36059), .B0(n28937), .Y(n28935)
         );
  NOR2BXL U19516 ( .AN(n36052), .B(conv_2[429]), .Y(n36055) );
  AOI2BB1XL U19517 ( .A0N(conv_2[427]), .A1N(n28904), .B0(n28906), .Y(n28923)
         );
  NOR2X1 U19518 ( .A(n28905), .B(n28910), .Y(n28924) );
  AOI2BB1XL U19519 ( .A0N(conv_2[426]), .A1N(n28929), .B0(n28906), .Y(n28904)
         );
  AOI2BB1XL U19520 ( .A0N(conv_2[425]), .A1N(n28893), .B0(n28906), .Y(n28929)
         );
  NOR2X1 U19521 ( .A(n28892), .B(n28891), .Y(n28930) );
  NOR2X1 U19522 ( .A(n35499), .B(n28125), .Y(n34488) );
  OR4XL U19523 ( .A(n34210), .B(conv_2[432]), .C(conv_2[431]), .D(n28906), .Y(
        n28911) );
  NOR2X1 U19524 ( .A(n33380), .B(n33321), .Y(n29486) );
  NOR2X1 U19525 ( .A(n33321), .B(n28076), .Y(n33377) );
  NOR2X1 U19526 ( .A(n34634), .B(n34635), .Y(n29531) );
  NOR2X1 U19527 ( .A(n33989), .B(n32016), .Y(n23212) );
  AOI2BB1XL U19528 ( .A0N(conv_2[382]), .A1N(n36023), .B0(n36025), .Y(n33673)
         );
  NOR2X1 U19529 ( .A(n34529), .B(n33675), .Y(n33672) );
  NOR2X1 U19530 ( .A(n34529), .B(n33417), .Y(n33414) );
  NOR2X1 U19531 ( .A(n29445), .B(n29449), .Y(n33417) );
  NOR2X1 U19532 ( .A(n33989), .B(n27532), .Y(n23988) );
  NOR2X1 U19533 ( .A(n29493), .B(n29492), .Y(n29495) );
  NOR2BXL U19534 ( .AN(n36018), .B(n36019), .Y(n24454) );
  OAI2BB1XL U19535 ( .A0N(n34568), .A1N(n34563), .B0(n34570), .Y(n36016) );
  NOR2BXL U19536 ( .AN(n36016), .B(conv_2[366]), .Y(n36019) );
  OAI2BB1XL U19537 ( .A0N(conv_2[365]), .A1N(n34564), .B0(n27273), .Y(n36018)
         );
  OR4XL U19538 ( .A(n34571), .B(conv_2[372]), .C(conv_2[371]), .D(n27273), .Y(
        n29467) );
  NOR2BXL U19539 ( .AN(n36011), .B(conv_2[356]), .Y(n36013) );
  AOI22XL U19540 ( .A0(n33925), .A1(n33924), .B0(n33931), .B1(n33926), .Y(
        n27993) );
  NOR2BXL U19541 ( .AN(n36004), .B(conv_2[341]), .Y(n36006) );
  OAI2BB1XL U19542 ( .A0N(conv_2[340]), .A1N(n29611), .B0(n35997), .Y(n36005)
         );
  NOR2BXL U19543 ( .AN(n35990), .B(n35991), .Y(n28102) );
  NOR2BXL U19544 ( .AN(n35989), .B(conv_2[336]), .Y(n35991) );
  OAI2BB1XL U19545 ( .A0N(conv_2[335]), .A1N(n28097), .B0(n35997), .Y(n35990)
         );
  OAI211X1 U19546 ( .A0(n23247), .A1(n34989), .B0(n22939), .C0(n22938), .Y(
        n34525) );
  AOI22XL U19547 ( .A0(n34827), .A1(n22937), .B0(n16755), .B1(n22936), .Y(
        n22939) );
  AOI2BB1XL U19548 ( .A0N(n35982), .A1N(n28064), .B0(n28063), .Y(n28060) );
  AOI2BB1XL U19549 ( .A0N(conv_2[320]), .A1N(n28050), .B0(n28051), .Y(n26352)
         );
  NAND2XL U19550 ( .A(n33979), .B(n28628), .Y(n35975) );
  NOR2BXL U19551 ( .AN(n35975), .B(conv_2[311]), .Y(n35978) );
  OAI2BB1XL U19552 ( .A0N(n28627), .A1N(conv_2[310]), .B0(n35970), .Y(n35977)
         );
  NAND2BXL U19553 ( .AN(conv_2[310]), .B(n19116), .Y(n28628) );
  OAI21XL U19554 ( .A0(conv_2[309]), .A1(n35968), .B0(n33979), .Y(n19116) );
  AOI2BB1XL U19555 ( .A0N(conv_2[306]), .A1N(n28917), .B0(n35970), .Y(n28898)
         );
  INVXL U19556 ( .A(n33979), .Y(n35970) );
  NOR2X1 U19557 ( .A(n19108), .B(n33989), .Y(n24181) );
  NAND2XL U19558 ( .A(n24181), .B(conv_2[300]), .Y(n24180) );
  NOR2BXL U19559 ( .AN(n35962), .B(conv_2[295]), .Y(n35965) );
  OAI2BB1XL U19560 ( .A0N(conv_2[294]), .A1N(n30979), .B0(n33135), .Y(n35964)
         );
  NOR2X1 U19561 ( .A(n30916), .B(n30917), .Y(n28093) );
  NOR2X1 U19562 ( .A(n30889), .B(n30892), .Y(n35956) );
  NAND2X1 U19563 ( .A(n22820), .B(n22819), .Y(n34455) );
  AOI22XL U19564 ( .A0(n26470), .A1(n22818), .B0(n28465), .B1(n22817), .Y(
        n22819) );
  AOI22XL U19565 ( .A0(n34827), .A1(n22850), .B0(n16755), .B1(n22849), .Y(
        n22820) );
  NOR2X1 U19566 ( .A(n28040), .B(n28039), .Y(n35949) );
  AOI2BB1XL U19567 ( .A0N(conv_2[278]), .A1N(n28033), .B0(n28883), .Y(n28038)
         );
  NAND2XL U19568 ( .A(n28739), .B(n34711), .Y(n28883) );
  AOI2BB1XL U19569 ( .A0N(conv_2[275]), .A1N(n28007), .B0(n28883), .Y(n18956)
         );
  AOI2BB1XL U19570 ( .A0N(n28011), .A1N(n28006), .B0(n35950), .Y(n28023) );
  NOR2X1 U19571 ( .A(n28189), .B(n28195), .Y(n28138) );
  NAND2XL U19572 ( .A(n28739), .B(n34422), .Y(n28161) );
  AOI21XL U19573 ( .A0(n28137), .A1(conv_2[262]), .B0(n28191), .Y(n28189) );
  NAND2BXL U19574 ( .AN(conv_2[262]), .B(n19046), .Y(n28190) );
  OR2XL U19575 ( .A(n28161), .B(n19044), .Y(n19046) );
  NOR2X1 U19576 ( .A(n33194), .B(n29455), .Y(n35940) );
  NOR2X1 U19577 ( .A(n33194), .B(n33199), .Y(n35941) );
  AOI2BB1XL U19578 ( .A0N(conv_2[245]), .A1N(n28258), .B0(n29455), .Y(n29143)
         );
  NOR2X1 U19579 ( .A(n29155), .B(n29159), .Y(n29598) );
  AOI2BB1XL U19580 ( .A0N(conv_2[231]), .A1N(n29173), .B0(n29174), .Y(n32875)
         );
  ADDFXL U19581 ( .A(conv_2[237]), .B(n32876), .CI(n31117), .CO(n33097), .S(
        n29600) );
  AOI21XL U19582 ( .A0(n30931), .A1(n30936), .B0(n30932), .Y(n31117) );
  AND2XL U19583 ( .A(n30437), .B(n35935), .Y(n35937) );
  OAI2BB1XL U19584 ( .A0N(conv_2[220]), .A1N(n30435), .B0(n31121), .Y(n35936)
         );
  NOR2X1 U19585 ( .A(n30430), .B(n31121), .Y(n30436) );
  NOR2X1 U19586 ( .A(n30429), .B(n30428), .Y(n30435) );
  NOR2X1 U19587 ( .A(n33770), .B(n33769), .Y(n33766) );
  AOI2BB1XL U19588 ( .A0N(conv_2[215]), .A1N(n29915), .B0(n29916), .Y(n29602)
         );
  NOR2X1 U19589 ( .A(n29916), .B(n29915), .Y(n29918) );
  NOR2X1 U19590 ( .A(n28660), .B(n23706), .Y(n34473) );
  ADDFXL U19591 ( .A(conv_2[206]), .B(n29935), .CI(n29921), .CO(n31310), .S(
        n29608) );
  AOI2BB1XL U19592 ( .A0N(conv_2[205]), .A1N(n29606), .B0(n29605), .Y(n29921)
         );
  AOI2BB1XL U19593 ( .A0N(conv_2[202]), .A1N(n29933), .B0(n35928), .Y(n35926)
         );
  AOI2BB1XL U19594 ( .A0N(conv_2[201]), .A1N(n35920), .B0(n35928), .Y(n29933)
         );
  NOR2X1 U19595 ( .A(n35921), .B(n35923), .Y(n29934) );
  AOI2BB1XL U19596 ( .A0N(conv_2[200]), .A1N(n29940), .B0(n35928), .Y(n35920)
         );
  NOR2X1 U19597 ( .A(n35928), .B(n27854), .Y(n29940) );
  AOI2BB1XL U19598 ( .A0N(conv_2[186]), .A1N(n29909), .B0(n30946), .Y(n29885)
         );
  AOI2BB1XL U19599 ( .A0N(conv_2[185]), .A1N(n29898), .B0(n30946), .Y(n29909)
         );
  NOR2X1 U19600 ( .A(n29897), .B(n29902), .Y(n29910) );
  AOI2BB1XL U19601 ( .A0N(conv_2[173]), .A1N(n29852), .B0(n29851), .Y(n30906)
         );
  NOR2X1 U19602 ( .A(n29851), .B(n29852), .Y(n29842) );
  NOR2X1 U19603 ( .A(n29831), .B(n29846), .Y(n29845) );
  AOI2BB1XL U19604 ( .A0N(conv_2[154]), .A1N(n23369), .B0(n23370), .Y(n24357)
         );
  NAND4X1 U19605 ( .A(n22176), .B(n22175), .C(n22174), .D(n22173), .Y(n34579)
         );
  AOI22XL U19606 ( .A0(n26470), .A1(n22936), .B0(n34827), .B1(n22305), .Y(
        n22174) );
  AOI22XL U19607 ( .A0(n28414), .A1(n22172), .B0(n35181), .B1(n22171), .Y(
        n22175) );
  NOR2X1 U19608 ( .A(n23296), .B(n23109), .Y(n34578) );
  NAND2XL U19609 ( .A(n35907), .B(n27973), .Y(n30082) );
  AOI2BB1XL U19610 ( .A0N(conv_2[144]), .A1N(n30087), .B0(n35899), .Y(n30094)
         );
  NOR2X1 U19611 ( .A(n30093), .B(n30088), .Y(n30095) );
  AOI2BB1XL U19612 ( .A0N(conv_2[143]), .A1N(n35905), .B0(n35899), .Y(n30087)
         );
  AOI2BB1XL U19613 ( .A0N(conv_2[142]), .A1N(n35897), .B0(n35899), .Y(n35905)
         );
  NOR2X1 U19614 ( .A(n35901), .B(n35898), .Y(n35906) );
  AOI2BB1XL U19615 ( .A0N(conv_2[141]), .A1N(n30076), .B0(n35899), .Y(n35897)
         );
  NAND2XL U19616 ( .A(n28739), .B(n34740), .Y(n35899) );
  NOR2X1 U19617 ( .A(n34426), .B(n34425), .Y(n34427) );
  AOI2BB1XL U19618 ( .A0N(conv_2[125]), .A1N(n34124), .B0(n30443), .Y(n33803)
         );
  NOR2X1 U19619 ( .A(n34344), .B(n33805), .Y(n33802) );
  NOR2X1 U19620 ( .A(n28948), .B(n23041), .Y(n34492) );
  ADDFXL U19621 ( .A(conv_2[132]), .B(n34344), .CI(n30067), .CO(n30444), .S(
        n24362) );
  AOI21XL U19622 ( .A0(n34355), .A1(n34350), .B0(n34351), .Y(n30067) );
  AOI2BB1XL U19623 ( .A0N(conv_2[111]), .A1N(n30143), .B0(n35884), .Y(n35882)
         );
  AOI2BB2XL U19624 ( .B0(n30210), .B1(n30225), .A0N(n30225), .A1N(n30206), .Y(
        n30216) );
  AOI32XL U19625 ( .A0(conv_2[99]), .A1(n30938), .A2(n30225), .B0(n30205), 
        .B1(n30938), .Y(n30212) );
  NAND2BXL U19626 ( .AN(conv_2[97]), .B(n19175), .Y(n30203) );
  OR2XL U19627 ( .A(n30225), .B(n19171), .Y(n28690) );
  NOR2X1 U19628 ( .A(n26509), .B(n19166), .Y(n34448) );
  AOI22XL U19629 ( .A0(n35130), .A1(n22123), .B0(n28465), .B1(n22803), .Y(
        n19163) );
  AOI22XL U19630 ( .A0(n16745), .A1(n22172), .B0(n35236), .B1(n22122), .Y(
        n19161) );
  AOI2BB1XL U19631 ( .A0N(conv_2[81]), .A1N(n35868), .B0(n30924), .Y(n30166)
         );
  AOI2BB1XL U19632 ( .A0N(conv_2[80]), .A1N(n30179), .B0(n30924), .Y(n35868)
         );
  NOR2X1 U19633 ( .A(n30240), .B(n30241), .Y(n30128) );
  NAND2XL U19634 ( .A(n31137), .B(n30162), .Y(n31135) );
  AOI2BB1XL U19635 ( .A0N(conv_2[51]), .A1N(n27819), .B0(n27820), .Y(n30872)
         );
  AOI2BB1XL U19636 ( .A0N(conv_2[36]), .A1N(n27728), .B0(n35862), .Y(n27711)
         );
  NOR2X1 U19637 ( .A(n33594), .B(n33596), .Y(n27729) );
  AND2XL U19638 ( .A(n33588), .B(n27707), .Y(n33592) );
  NOR2X1 U19639 ( .A(n33588), .B(n27707), .Y(n33594) );
  NOR2X1 U19640 ( .A(conv_2[26]), .B(n27837), .Y(n27843) );
  NOR2X1 U19641 ( .A(n27843), .B(n27836), .Y(n27842) );
  OR2XL U19642 ( .A(n33620), .B(n27555), .Y(n29075) );
  NOR2X1 U19643 ( .A(n30195), .B(n33989), .Y(n24199) );
  NOR2X1 U19644 ( .A(n28783), .B(n28779), .Y(n28785) );
  NOR2X1 U19645 ( .A(n33569), .B(n29583), .Y(n28778) );
  NOR2X1 U19646 ( .A(n29587), .B(n29582), .Y(n33570) );
  INVXL U19647 ( .A(n29583), .Y(n33571) );
  NAND2XL U19648 ( .A(n27691), .B(n28739), .Y(n29583) );
  NOR2X1 U19649 ( .A(n33989), .B(n35857), .Y(n24004) );
  NAND2X1 U19650 ( .A(n22896), .B(filter_2_bias[0]), .Y(n34583) );
  NOR2X1 U19651 ( .A(n27568), .B(n28959), .Y(n33716) );
  NOR4BXL U19652 ( .AN(n21122), .B(n21121), .C(n21120), .D(n21119), .Y(n21457)
         );
  OAI21XL U19653 ( .A0(n35229), .A1(n21455), .B0(n35227), .Y(n35014) );
  AOI222XL U19654 ( .A0(n21454), .A1(n21453), .B0(n21454), .B1(n21452), .C0(
        n21453), .C1(n21451), .Y(n21455) );
  INVXL U19655 ( .A(n34921), .Y(n25853) );
  OAI21XL U19656 ( .A0(n35229), .A1(n19606), .B0(n35227), .Y(n35026) );
  AOI222XL U19657 ( .A0(n19605), .A1(n19604), .B0(n19605), .B1(n19603), .C0(
        n19604), .C1(n19602), .Y(n19606) );
  AOI211XL U19658 ( .A0(n34963), .A1(n34986), .B0(n26161), .C0(n26160), .Y(
        n26296) );
  OAI21XL U19659 ( .A0(n35229), .A1(n26294), .B0(n35227), .Y(n34945) );
  AOI222XL U19660 ( .A0(n26293), .A1(n26292), .B0(n26293), .B1(n26291), .C0(
        n26292), .C1(n26290), .Y(n26294) );
  OAI21XL U19661 ( .A0(n35229), .A1(n18722), .B0(n35227), .Y(n24569) );
  AOI222XL U19662 ( .A0(n18721), .A1(n18720), .B0(n18721), .B1(n18719), .C0(
        n18720), .C1(n18718), .Y(n18722) );
  OR2XL U19663 ( .A(n28296), .B(n28295), .Y(n35003) );
  OAI2BB1XL U19664 ( .A0N(n28391), .A1N(n28390), .B0(n35227), .Y(n35010) );
  AOI222XL U19665 ( .A0(n28389), .A1(n28388), .B0(n28389), .B1(n28387), .C0(
        n28388), .C1(n28386), .Y(n28390) );
  AOI211XL U19666 ( .A0(n34827), .A1(n35175), .B0(n28269), .C0(n28268), .Y(
        n28389) );
  INVXL U19667 ( .A(n35010), .Y(n35006) );
  AOI211XL U19668 ( .A0(n26470), .A1(n25691), .B0(n25690), .C0(n25689), .Y(
        n25811) );
  OAI21XL U19669 ( .A0(n35229), .A1(n25809), .B0(n35227), .Y(n35022) );
  INVXL U19670 ( .A(n33429), .Y(n34498) );
  NOR2X1 U19671 ( .A(n33429), .B(n23545), .Y(n28620) );
  AOI2BB1XL U19672 ( .A0N(conv_3[514]), .A1N(n24459), .B0(n24458), .Y(n24478)
         );
  NAND2XL U19673 ( .A(n35838), .B(n33856), .Y(n33919) );
  AOI2BB1XL U19674 ( .A0N(conv_3[503]), .A1N(n32082), .B0(n33918), .Y(n32076)
         );
  AOI2BB1XL U19675 ( .A0N(conv_3[501]), .A1N(n35836), .B0(n33918), .Y(n27629)
         );
  NAND2XL U19676 ( .A(n31924), .B(n33424), .Y(n33918) );
  AOI2BB1XL U19677 ( .A0N(conv_3[500]), .A1N(n32071), .B0(n33918), .Y(n35836)
         );
  NOR2X1 U19678 ( .A(n32070), .B(n32075), .Y(n35837) );
  NOR2X1 U19679 ( .A(n27620), .B(n33422), .Y(n31381) );
  NOR2X1 U19680 ( .A(n31549), .B(n31548), .Y(n35830) );
  AOI2BB1XL U19681 ( .A0N(conv_3[484]), .A1N(n23773), .B0(n23772), .Y(n27614)
         );
  NOR2X1 U19682 ( .A(n35810), .B(n32185), .Y(n19027) );
  AOI2BB1XL U19683 ( .A0N(conv_3[472]), .A1N(n32333), .B0(n32334), .Y(n33011)
         );
  NOR2X1 U19684 ( .A(n31517), .B(n19062), .Y(n35795) );
  OAI211X1 U19685 ( .A0(n22800), .A1(n34989), .B0(n19057), .C0(n19056), .Y(
        n34444) );
  AOI21XL U19686 ( .A0(n16755), .A1(n22804), .B0(n19055), .Y(n19056) );
  OAI211XL U19687 ( .A0(n22807), .A1(n16701), .B0(n19054), .C0(n19053), .Y(
        n19055) );
  NOR2X1 U19688 ( .A(conv_3[446]), .B(n31950), .Y(n31945) );
  NOR2X1 U19689 ( .A(n31945), .B(n31949), .Y(n31943) );
  OAI211X1 U19690 ( .A0(n22892), .A1(n35135), .B0(n22891), .C0(n22890), .Y(
        n34224) );
  NOR3XL U19691 ( .A(n32158), .B(conv_3[432]), .C(n35775), .Y(n32590) );
  AOI2BB1XL U19692 ( .A0N(conv_3[428]), .A1N(n31701), .B0(n35775), .Y(n35773)
         );
  AOI2BB1XL U19693 ( .A0N(conv_3[427]), .A1N(n35767), .B0(n35775), .Y(n31701)
         );
  NOR2X1 U19694 ( .A(n35770), .B(n35768), .Y(n31702) );
  AOI2BB1XL U19695 ( .A0N(conv_3[425]), .A1N(n32576), .B0(n35775), .Y(n33786)
         );
  NOR2X1 U19696 ( .A(n33790), .B(n33789), .Y(n33785) );
  NOR2X1 U19697 ( .A(n32575), .B(n32579), .Y(n33789) );
  NOR2X1 U19698 ( .A(conv_3[433]), .B(n32590), .Y(n32589) );
  OR2XL U19699 ( .A(n32558), .B(n31994), .Y(n31999) );
  INVXL U19700 ( .A(n28070), .Y(n34229) );
  OR2XL U19701 ( .A(n33695), .B(n33222), .Y(n33697) );
  NOR2X1 U19702 ( .A(n33222), .B(n33221), .Y(n33696) );
  NOR2X1 U19703 ( .A(n32037), .B(n32038), .Y(n32034) );
  NAND3BX1 U19704 ( .AN(n23020), .B(n23019), .C(n23018), .Y(n27990) );
  AOI22XL U19705 ( .A0(n23055), .A1(n23277), .B0(n23017), .B1(n23273), .Y(
        n23018) );
  AOI22XL U19706 ( .A0(n25766), .A1(n23275), .B0(n34906), .B1(n23782), .Y(
        n23019) );
  OAI22XL U19707 ( .A0(n23282), .A1(n25853), .B0(N18471), .B1(n23285), .Y(
        n23020) );
  NOR2X1 U19708 ( .A(n32197), .B(n32198), .Y(n31388) );
  AND2XL U19709 ( .A(n31386), .B(n31385), .Y(n32525) );
  NOR2X1 U19710 ( .A(n31691), .B(n27532), .Y(n23070) );
  AOI2BB1XL U19711 ( .A0N(conv_3[378]), .A1N(n24202), .B0(n24203), .Y(n23069)
         );
  NOR2X1 U19712 ( .A(n27532), .B(n27531), .Y(n27533) );
  NOR2X1 U19713 ( .A(conv_3[371]), .B(n31631), .Y(n31644) );
  AOI2BB1XL U19714 ( .A0N(conv_3[366]), .A1N(n31660), .B0(n35761), .Y(n31654)
         );
  NAND2XL U19715 ( .A(conv_3[360]), .B(n31330), .Y(n31329) );
  AOI2BB1XL U19716 ( .A0N(conv_3[352]), .A1N(n31466), .B0(n32130), .Y(n33749)
         );
  NOR2X1 U19717 ( .A(conv_3[353]), .B(n33749), .Y(n33750) );
  NOR2X1 U19718 ( .A(n31468), .B(n31467), .Y(n33751) );
  AOI2BB1XL U19719 ( .A0N(conv_3[351]), .A1N(n31450), .B0(n32130), .Y(n31466)
         );
  NAND2XL U19720 ( .A(n31924), .B(n34762), .Y(n32130) );
  NOR2X1 U19721 ( .A(n27620), .B(n26717), .Y(n27043) );
  NAND2XL U19722 ( .A(n31980), .B(n31970), .Y(n31982) );
  OAI2BB1XL U19723 ( .A0N(conv_3[340]), .A1N(n31975), .B0(n31967), .Y(n31981)
         );
  AOI2BB1XL U19724 ( .A0N(n31980), .A1N(n31975), .B0(n31974), .Y(n31977) );
  NOR2X1 U19725 ( .A(n31967), .B(n23769), .Y(n35746) );
  NOR2X1 U19726 ( .A(n27620), .B(n34522), .Y(n30615) );
  NOR2BXL U19727 ( .AN(n33280), .B(n31919), .Y(n31921) );
  ADDFXL U19728 ( .A(conv_3[324]), .B(n33842), .CI(n32528), .CO(n31915), .S(
        n32529) );
  AOI2BB1XL U19729 ( .A0N(n35739), .A1N(conv_3[323]), .B0(n35740), .Y(n32528)
         );
  NOR2X1 U19730 ( .A(n31907), .B(n33281), .Y(n33839) );
  NOR2X1 U19731 ( .A(n33842), .B(n33841), .Y(n33838) );
  ADDFXL U19732 ( .A(conv_3[310]), .B(n35732), .CI(n32613), .CO(n32609), .S(
        n32615) );
  AOI21XL U19733 ( .A0(n32540), .A1(n32535), .B0(n32536), .Y(n32613) );
  NOR2X1 U19734 ( .A(n35732), .B(n35733), .Y(n35731) );
  ADDFXL U19735 ( .A(conv_3[306]), .B(n35732), .CI(n32549), .CO(n35733), .S(
        n32550) );
  AOI2BB1XL U19736 ( .A0N(conv_3[305]), .A1N(n31443), .B0(n31444), .Y(n32549)
         );
  NOR2X1 U19737 ( .A(n19108), .B(n23216), .Y(n27058) );
  ADDFXL U19738 ( .A(conv_3[289]), .B(n31873), .CI(n31872), .CO(n31888), .S(
        n23067) );
  NOR2X1 U19739 ( .A(n31691), .B(n31871), .Y(n31873) );
  AOI2BB1XL U19740 ( .A0N(conv_3[288]), .A1N(n23666), .B0(n23667), .Y(n31872)
         );
  NOR2X1 U19741 ( .A(n35720), .B(n31888), .Y(n31877) );
  OR4XL U19742 ( .A(n34479), .B(conv_3[296]), .C(conv_3[297]), .D(n31896), .Y(
        n32235) );
  NOR2X1 U19743 ( .A(n32618), .B(n31757), .Y(n31756) );
  ADDFXL U19744 ( .A(conv_3[279]), .B(n32618), .CI(n32617), .CO(n31757), .S(
        n32620) );
  AOI2BB1XL U19745 ( .A0N(conv_3[278]), .A1N(n31738), .B0(n31739), .Y(n32617)
         );
  NOR2X1 U19746 ( .A(n33994), .B(n22858), .Y(n34710) );
  NOR2XL U19747 ( .A(n33480), .B(n33481), .Y(n33227) );
  NOR2BXL U19748 ( .AN(n35712), .B(conv_3[265]), .Y(n35715) );
  NOR2X1 U19749 ( .A(n32101), .B(n32100), .Y(n33006) );
  AOI2BB1XL U19750 ( .A0N(conv_3[262]), .A1N(n29106), .B0(n33478), .Y(n28726)
         );
  NOR2X1 U19751 ( .A(conv_3[263]), .B(n28726), .Y(n32102) );
  AOI2BB1XL U19752 ( .A0N(conv_3[261]), .A1N(n29130), .B0(n33478), .Y(n29106)
         );
  NOR2X1 U19753 ( .A(n29131), .B(n29135), .Y(n29107) );
  AOI2BB1XL U19754 ( .A0N(conv_3[260]), .A1N(n29112), .B0(n33478), .Y(n29130)
         );
  NOR2X1 U19755 ( .A(n33478), .B(n28724), .Y(n29112) );
  NOR2X1 U19756 ( .A(n27620), .B(n28721), .Y(n30607) );
  NOR2X1 U19757 ( .A(conv_3[251]), .B(n35705), .Y(n35709) );
  NOR2X1 U19758 ( .A(n35702), .B(n35699), .Y(n29118) );
  AOI2BB1XL U19759 ( .A0N(conv_3[249]), .A1N(n35698), .B0(n35700), .Y(n28800)
         );
  NOR2X1 U19760 ( .A(n35693), .B(n29118), .Y(n28799) );
  AOI2BB1XL U19761 ( .A0N(conv_3[248]), .A1N(n35691), .B0(n35700), .Y(n35698)
         );
  AOI2BB1XL U19762 ( .A0N(conv_3[247]), .A1N(n35685), .B0(n35700), .Y(n35691)
         );
  NOR2X1 U19763 ( .A(n35688), .B(n35686), .Y(n35692) );
  AOI2BB1XL U19764 ( .A0N(conv_3[246]), .A1N(n35679), .B0(n35700), .Y(n35685)
         );
  NAND2XL U19765 ( .A(n31924), .B(n33535), .Y(n35700) );
  AOI2BB1XL U19766 ( .A0N(conv_3[245]), .A1N(n34246), .B0(n35700), .Y(n35679)
         );
  NOR2X1 U19767 ( .A(n34245), .B(n34249), .Y(n35680) );
  NOR2X1 U19768 ( .A(n27620), .B(n24021), .Y(n30603) );
  NAND2XL U19769 ( .A(n35673), .B(n33316), .Y(n33879) );
  AOI2BB1XL U19770 ( .A0N(conv_3[234]), .A1N(n30689), .B0(n33878), .Y(n31060)
         );
  NOR2X1 U19771 ( .A(n30694), .B(n30690), .Y(n31061) );
  AOI2BB1XL U19772 ( .A0N(conv_3[233]), .A1N(n35671), .B0(n33878), .Y(n30689)
         );
  AOI2BB1XL U19773 ( .A0N(conv_3[232]), .A1N(n32094), .B0(n33878), .Y(n35671)
         );
  AOI2BB1XL U19774 ( .A0N(conv_3[231]), .A1N(n32088), .B0(n33878), .Y(n32094)
         );
  NAND2XL U19775 ( .A(n34461), .B(n31924), .Y(n33878) );
  AOI2BB1XL U19776 ( .A0N(conv_3[230]), .A1N(n29162), .B0(n33878), .Y(n32088)
         );
  NOR2X1 U19777 ( .A(n29161), .B(n29160), .Y(n32089) );
  NOR2X1 U19778 ( .A(n32058), .B(n34649), .Y(n31536) );
  NOR2X1 U19779 ( .A(n28660), .B(n23617), .Y(n27492) );
  NAND2XL U19780 ( .A(n35653), .B(n31850), .Y(n31860) );
  NOR2X1 U19781 ( .A(n31849), .B(n31848), .Y(n35651) );
  NOR2X1 U19782 ( .A(n31847), .B(n31846), .Y(n35652) );
  NOR2X1 U19783 ( .A(n31866), .B(n31865), .Y(n31868) );
  NOR2X1 U19784 ( .A(n27848), .B(n27620), .Y(n30842) );
  NAND2XL U19785 ( .A(n31591), .B(conv_3[188]), .Y(n31609) );
  NOR2X1 U19786 ( .A(n31596), .B(n31601), .Y(n31591) );
  AOI2BB1XL U19787 ( .A0N(conv_3[185]), .A1N(n31614), .B0(n31615), .Y(n32648)
         );
  NOR3XL U19788 ( .A(n32222), .B(conv_3[177]), .C(n32221), .Y(n32644) );
  NOR2X1 U19789 ( .A(n31579), .B(n31578), .Y(n32220) );
  NOR2X1 U19790 ( .A(n31577), .B(n31578), .Y(n31570) );
  AOI2BB1XL U19791 ( .A0N(conv_3[174]), .A1N(n31573), .B0(n32221), .Y(n35637)
         );
  NOR2X1 U19792 ( .A(n35636), .B(n35635), .Y(n35638) );
  ADDFXL U19793 ( .A(conv_3[173]), .B(n35639), .CI(n32658), .CO(n31573), .S(
        n32659) );
  NOR2BXL U19794 ( .AN(n35631), .B(n35632), .Y(n32658) );
  INVX2 U19795 ( .A(n36056), .Y(n36001) );
  NOR2X1 U19796 ( .A(n32314), .B(n32320), .Y(n32291) );
  AOI21XL U19797 ( .A0(conv_3[160]), .A1(n32303), .B0(n32316), .Y(n32314) );
  OR2XL U19798 ( .A(n32252), .B(n32251), .Y(n32302) );
  NOR2X1 U19799 ( .A(n32251), .B(n32296), .Y(n32303) );
  AOI2BB1XL U19800 ( .A0N(conv_3[156]), .A1N(n32308), .B0(n32252), .Y(n29749)
         );
  NAND2XL U19801 ( .A(n31924), .B(n34579), .Y(n32252) );
  AOI2BB1XL U19802 ( .A0N(conv_3[155]), .A1N(n32285), .B0(n32252), .Y(n32308)
         );
  NOR2X1 U19803 ( .A(n32284), .B(n32289), .Y(n32309) );
  NOR2X1 U19804 ( .A(conv_3[146]), .B(n33967), .Y(n32788) );
  AOI2BB1XL U19805 ( .A0N(conv_3[141]), .A1N(n31713), .B0(n31714), .Y(n28623)
         );
  NOR2X1 U19806 ( .A(n35622), .B(n35623), .Y(n35621) );
  NAND2XL U19807 ( .A(n30838), .B(conv_3[120]), .Y(n30837) );
  AOI2BB1XL U19808 ( .A0N(conv_3[111]), .A1N(n31784), .B0(n31786), .Y(n31797)
         );
  AOI2BB1XL U19809 ( .A0N(conv_3[110]), .A1N(n31774), .B0(n31786), .Y(n31784)
         );
  INVXL U19810 ( .A(n34196), .Y(n31786) );
  NOR2X1 U19811 ( .A(n31786), .B(n31769), .Y(n31774) );
  NOR2X1 U19812 ( .A(n27620), .B(n34715), .Y(n30830) );
  NAND2XL U19813 ( .A(n30830), .B(conv_3[105]), .Y(n30829) );
  NOR2X1 U19814 ( .A(n33742), .B(n35615), .Y(n31673) );
  NOR2X1 U19815 ( .A(n34186), .B(n33743), .Y(n33740) );
  NOR2X1 U19816 ( .A(n26509), .B(n27620), .Y(n30834) );
  NAND2X1 U19817 ( .A(n30834), .B(conv_3[90]), .Y(n30833) );
  NAND2XL U19818 ( .A(n31842), .B(n31829), .Y(n31840) );
  AOI2BB1XL U19819 ( .A0N(conv_3[84]), .A1N(n35605), .B0(n35607), .Y(n31816)
         );
  AOI2BB1XL U19820 ( .A0N(conv_3[83]), .A1N(n31810), .B0(n35607), .Y(n35605)
         );
  AOI2BB1XL U19821 ( .A0N(conv_3[81]), .A1N(n31821), .B0(n35607), .Y(n31833)
         );
  NAND2XL U19822 ( .A(n31924), .B(n34438), .Y(n35607) );
  INVX2 U19823 ( .A(n34438), .Y(n33020) );
  NOR2XL U19824 ( .A(n35599), .B(n32164), .Y(n31421) );
  NAND2XL U19825 ( .A(conv_3[67]), .B(n35601), .Y(n31491) );
  ADDFXL U19826 ( .A(conv_3[66]), .B(n35599), .CI(n32542), .CO(n35600), .S(
        n32543) );
  ADDFXL U19827 ( .A(conv_3[65]), .B(n35599), .CI(n32605), .CO(n32542), .S(
        n32607) );
  AOI2BB1XL U19828 ( .A0N(conv_3[64]), .A1N(n31420), .B0(n31419), .Y(n32605)
         );
  INVXL U19829 ( .A(n31418), .Y(n34699) );
  NOR2XL U19830 ( .A(n31418), .B(n23895), .Y(n34698) );
  NOR2X1 U19831 ( .A(n32179), .B(n32178), .Y(n33820) );
  NOR2X1 U19832 ( .A(n33824), .B(n33823), .Y(n33819) );
  INVXL U19833 ( .A(n34507), .Y(n27799) );
  NOR2X1 U19834 ( .A(n33449), .B(n31239), .Y(n31238) );
  ADDFXL U19835 ( .A(conv_3[41]), .B(n33449), .CI(n31222), .CO(n31239), .S(
        n24471) );
  AOI2BB1XL U19836 ( .A0N(conv_3[40]), .A1N(n31232), .B0(n31233), .Y(n31222)
         );
  NOR2X1 U19837 ( .A(conv_3[37]), .B(n33446), .Y(n33447) );
  NOR2X1 U19838 ( .A(n31245), .B(n31249), .Y(n33448) );
  AOI2BB1XL U19839 ( .A0N(conv_3[36]), .A1N(n31244), .B0(n35591), .Y(n33446)
         );
  NOR2X1 U19840 ( .A(n33449), .B(n33448), .Y(n33445) );
  NOR2X1 U19841 ( .A(n35585), .B(n35591), .Y(n31244) );
  NOR2X1 U19842 ( .A(n35591), .B(n24470), .Y(n35582) );
  NOR2X1 U19843 ( .A(n31251), .B(n31250), .Y(n31257) );
  NOR2X1 U19844 ( .A(n31262), .B(n31266), .Y(n31268) );
  AOI2BB1XL U19845 ( .A0N(conv_3[19]), .A1N(n30197), .B0(n30196), .Y(n33001)
         );
  AOI22XL U19846 ( .A0(n16745), .A1(n22399), .B0(n26263), .B1(n22845), .Y(
        n21105) );
  AOI211XL U19847 ( .A0(n35181), .A1(n22397), .B0(n21097), .C0(n21096), .Y(
        n21104) );
  AOI22XL U19848 ( .A0(n35130), .A1(n22848), .B0(n28465), .B1(n22849), .Y(
        n21103) );
  AOI222XL U19849 ( .A0(conv_3[8]), .A1(n34379), .B0(n32996), .B1(n24372), 
        .C0(n31196), .C1(n31194), .Y(n31159) );
  ADDFXL U19850 ( .A(conv_3[4]), .B(n24369), .CI(n24368), .CO(n28687), .S(
        n23757) );
  NOR2X1 U19851 ( .A(n31691), .B(n35857), .Y(n24369) );
  NAND2XL U19852 ( .A(conv_3[0]), .B(n31027), .Y(n31026) );
  NAND2X1 U19853 ( .A(n22896), .B(filter_3_bias[0]), .Y(n34755) );
  INVXL U19854 ( .A(n36114), .Y(n20180) );
  INVX2 U19855 ( .A(n30392), .Y(n36107) );
  OAI2BB1XL U19856 ( .A0N(n20168), .A1N(n20167), .B0(n20166), .Y(n36139) );
  OAI21XL U19857 ( .A0(n20179), .A1(in_data[10]), .B0(n20178), .Y(n36142) );
  OAI2BB1XL U19858 ( .A0N(n20178), .A1N(n20172), .B0(n20171), .Y(n36145) );
  OAI21XL U19859 ( .A0(n20170), .A1(in_data[12]), .B0(n20174), .Y(n36148) );
  XOR2XL U19860 ( .A(in_data[13]), .B(n20174), .Y(n36151) );
  NOR2X1 U19861 ( .A(n35261), .B(n35260), .Y(n35264) );
  OAI21XL U19862 ( .A0(n35259), .A1(n36042), .B0(n35261), .Y(n35267) );
  NOR2X1 U19863 ( .A(in_data[3]), .B(in_data[4]), .Y(n25083) );
  NOR3XL U19864 ( .A(n18174), .B(n18175), .C(n18173), .Y(n18181) );
  OAI21XL U19865 ( .A0(n18177), .A1(n18176), .B0(cs[1]), .Y(n18178) );
  NAND2XL U19866 ( .A(n18773), .B(n26850), .Y(n18167) );
  INVXL U19867 ( .A(n19245), .Y(n19229) );
  OAI31XL U19868 ( .A0(n19226), .A1(n19225), .A2(n19224), .B0(n19223), .Y(
        n16641) );
  AOI22XL U19869 ( .A0(N29498), .A1(n35256), .B0(n19222), .B1(n19221), .Y(
        n19223) );
  AOI211XL U19870 ( .A0(n19247), .A1(n18172), .B0(n20358), .C0(n19242), .Y(
        N30142) );
  NAND2XL U19871 ( .A(n33078), .B(n33077), .Y(n16504) );
  OAI2BB2XL U19872 ( .B0(n33074), .B1(n33073), .A0N(n33074), .A1N(n33073), .Y(
        n33076) );
  AOI22XL U19873 ( .A0(n33563), .A1(n33562), .B0(affine_1[19]), .B1(n33561), 
        .Y(n33565) );
  OAI22XL U19874 ( .A0(n16645), .A1(n32962), .B0(n32961), .B1(n26853), .Y(
        n14106) );
  OAI22XL U19875 ( .A0(n16650), .A1(n32961), .B0(n32960), .B1(n26853), .Y(
        n14107) );
  OAI22XL U19876 ( .A0(n16645), .A1(n32960), .B0(n32958), .B1(n26853), .Y(
        n14108) );
  OAI22XL U19877 ( .A0(n32967), .A1(n32958), .B0(n32957), .B1(n26853), .Y(
        n14109) );
  OAI22XL U19878 ( .A0(n16645), .A1(n32957), .B0(n32955), .B1(n26853), .Y(
        n14110) );
  OAI22XL U19879 ( .A0(n31084), .A1(n32955), .B0(n32954), .B1(n26853), .Y(
        n14111) );
  OAI22XL U19880 ( .A0(n32491), .A1(n32954), .B0(n32953), .B1(n26853), .Y(
        n14112) );
  OAI22XL U19881 ( .A0(n31071), .A1(n32953), .B0(n32952), .B1(n26853), .Y(
        n14113) );
  OAI22XL U19882 ( .A0(n16650), .A1(n32952), .B0(n32951), .B1(n26853), .Y(
        n14114) );
  OAI22XL U19883 ( .A0(n26906), .A1(n32951), .B0(n32950), .B1(n26853), .Y(
        n14115) );
  OAI22XL U19884 ( .A0(n16645), .A1(n32950), .B0(n32947), .B1(n26853), .Y(
        n14116) );
  OAI22XL U19885 ( .A0(n31077), .A1(n32947), .B0(n32944), .B1(n26853), .Y(
        n14117) );
  OAI22XL U19886 ( .A0(n16650), .A1(n32944), .B0(n32943), .B1(n26853), .Y(
        n14118) );
  OAI22XL U19887 ( .A0(n32491), .A1(n32943), .B0(n32942), .B1(n26853), .Y(
        n14119) );
  OAI22XL U19888 ( .A0(n16650), .A1(n32942), .B0(n32941), .B1(n26853), .Y(
        n14120) );
  OAI22XL U19889 ( .A0(n31084), .A1(n32941), .B0(n32937), .B1(n26853), .Y(
        n14121) );
  OAI22XL U19890 ( .A0(n32491), .A1(n32937), .B0(n32936), .B1(n26853), .Y(
        n14122) );
  OAI22XL U19891 ( .A0(n16645), .A1(n32936), .B0(n32935), .B1(n26853), .Y(
        n14123) );
  OAI22XL U19892 ( .A0(n31071), .A1(n32935), .B0(n32934), .B1(n26853), .Y(
        n14124) );
  OAI22XL U19893 ( .A0(n31071), .A1(n32934), .B0(n32933), .B1(n26853), .Y(
        n14125) );
  OAI22XL U19894 ( .A0(n31071), .A1(n32933), .B0(n32932), .B1(n26853), .Y(
        n14126) );
  OAI22XL U19895 ( .A0(n16645), .A1(n32932), .B0(n32931), .B1(n26853), .Y(
        n14127) );
  OAI22XL U19896 ( .A0(n32967), .A1(n32931), .B0(n32928), .B1(n26853), .Y(
        n14128) );
  OAI22XL U19897 ( .A0(n16645), .A1(n32928), .B0(n32927), .B1(n26853), .Y(
        n14129) );
  OAI22XL U19898 ( .A0(n16650), .A1(n32927), .B0(n32926), .B1(n26853), .Y(
        n14130) );
  OAI22XL U19899 ( .A0(n16650), .A1(n32926), .B0(n32925), .B1(n26853), .Y(
        n14131) );
  OAI22XL U19900 ( .A0(n16645), .A1(n32925), .B0(n32924), .B1(n26853), .Y(
        n14132) );
  OAI22XL U19901 ( .A0(n32967), .A1(n32924), .B0(n32964), .B1(n26853), .Y(
        n14133) );
  OAI22XL U19902 ( .A0(n16645), .A1(n32964), .B0(n32963), .B1(n26853), .Y(
        n14134) );
  OAI22XL U19903 ( .A0(n26906), .A1(n32963), .B0(n32920), .B1(n26853), .Y(
        n14135) );
  OAI22XL U19904 ( .A0(n16650), .A1(n32920), .B0(n32919), .B1(n26853), .Y(
        n14136) );
  OAI22XL U19905 ( .A0(n16645), .A1(n32919), .B0(n32915), .B1(n26853), .Y(
        n14137) );
  OAI22XL U19906 ( .A0(n32967), .A1(n32915), .B0(n32914), .B1(n26853), .Y(
        n14138) );
  OAI22XL U19907 ( .A0(n31077), .A1(n32914), .B0(n32913), .B1(n26853), .Y(
        n14139) );
  OAI22XL U19908 ( .A0(n16650), .A1(n32913), .B0(n32912), .B1(n26853), .Y(
        n14140) );
  OAI22XL U19909 ( .A0(n16650), .A1(n32909), .B0(n32949), .B1(n26853), .Y(
        n14159) );
  OAI22XL U19910 ( .A0(n16645), .A1(n32949), .B0(n32948), .B1(n26853), .Y(
        n14160) );
  OAI22XL U19911 ( .A0(n32967), .A1(n32948), .B0(n32946), .B1(n26853), .Y(
        n14161) );
  OAI22XL U19912 ( .A0(n16645), .A1(n32946), .B0(n32945), .B1(n26853), .Y(
        n14162) );
  OAI22XL U19913 ( .A0(n31071), .A1(n32945), .B0(n32904), .B1(n26853), .Y(
        n14163) );
  OAI22XL U19914 ( .A0(n16645), .A1(n32904), .B0(n32903), .B1(n26853), .Y(
        n14164) );
  OAI22XL U19915 ( .A0(n16645), .A1(n32903), .B0(n32940), .B1(n26853), .Y(
        n14165) );
  OAI22XL U19916 ( .A0(n32967), .A1(n32940), .B0(n32939), .B1(n26853), .Y(
        n14166) );
  OAI22XL U19917 ( .A0(n16650), .A1(n32939), .B0(n32938), .B1(n26853), .Y(
        n14167) );
  OAI22XL U19918 ( .A0(n32491), .A1(n32938), .B0(n32900), .B1(n26853), .Y(
        n14168) );
  OAI22XL U19919 ( .A0(n32967), .A1(n32900), .B0(n32899), .B1(n26853), .Y(
        n14169) );
  OAI22XL U19920 ( .A0(n16650), .A1(n32899), .B0(n32896), .B1(n26853), .Y(
        n14170) );
  OAI22XL U19921 ( .A0(n16650), .A1(n32896), .B0(n32895), .B1(n26853), .Y(
        n14171) );
  OAI22XL U19922 ( .A0(n31084), .A1(n32895), .B0(n32908), .B1(n26853), .Y(
        n14172) );
  OAI22XL U19923 ( .A0(n16645), .A1(n32908), .B0(n32907), .B1(n26853), .Y(
        n14173) );
  OAI22XL U19924 ( .A0(n16645), .A1(n32907), .B0(n32916), .B1(n26853), .Y(
        n14174) );
  OAI22XL U19925 ( .A0(n16645), .A1(n32916), .B0(n32918), .B1(n26853), .Y(
        n14175) );
  OAI22XL U19926 ( .A0(n16645), .A1(n32918), .B0(n32917), .B1(n26853), .Y(
        n14176) );
  OAI22XL U19927 ( .A0(n16645), .A1(n32917), .B0(n32921), .B1(n26853), .Y(
        n14177) );
  OAI22XL U19928 ( .A0(n32491), .A1(n32921), .B0(n32923), .B1(n26853), .Y(
        n14178) );
  OAI22XL U19929 ( .A0(n16645), .A1(n32923), .B0(n32922), .B1(n26853), .Y(
        n14179) );
  OAI22XL U19930 ( .A0(n31084), .A1(n32922), .B0(n32902), .B1(n26853), .Y(
        n14180) );
  OAI22XL U19931 ( .A0(n31071), .A1(n32902), .B0(n32901), .B1(n26853), .Y(
        n14181) );
  OAI22XL U19932 ( .A0(n16645), .A1(n32901), .B0(n32906), .B1(n26853), .Y(
        n14182) );
  OAI22XL U19933 ( .A0(n16645), .A1(n32906), .B0(n32905), .B1(n26853), .Y(
        n14183) );
  OAI22XL U19934 ( .A0(n32967), .A1(n32905), .B0(n32930), .B1(n26853), .Y(
        n14184) );
  OAI22XL U19935 ( .A0(n32967), .A1(n32930), .B0(n32929), .B1(n26853), .Y(
        n14185) );
  OAI22XL U19936 ( .A0(n32967), .A1(n32929), .B0(n36151), .B1(n26853), .Y(
        n14186) );
  OAI22XL U19937 ( .A0(n32967), .A1(n32910), .B0(n32966), .B1(n26853), .Y(
        n14187) );
  OAI22XL U19938 ( .A0(n32967), .A1(n32966), .B0(n32965), .B1(n26853), .Y(
        n14188) );
  OAI22XL U19939 ( .A0(n32967), .A1(n32965), .B0(n32911), .B1(n26853), .Y(
        n14189) );
  OAI22XL U19940 ( .A0(n32967), .A1(n32911), .B0(n32898), .B1(n26853), .Y(
        n14190) );
  OAI22XL U19941 ( .A0(n32967), .A1(n32898), .B0(n32897), .B1(n26853), .Y(
        n14191) );
  OAI22XL U19942 ( .A0(n16645), .A1(n32956), .B0(n32959), .B1(n26853), .Y(
        n14218) );
  OAI22XL U19943 ( .A0(n31077), .A1(n32959), .B0(n32973), .B1(n26853), .Y(
        n14219) );
  OAI22XL U19944 ( .A0(n16645), .A1(n32973), .B0(n32972), .B1(n26853), .Y(
        n14220) );
  OAI22XL U19945 ( .A0(n16645), .A1(n32972), .B0(n32975), .B1(n26853), .Y(
        n14221) );
  OAI22XL U19946 ( .A0(n16645), .A1(n32975), .B0(n32974), .B1(n26853), .Y(
        n14222) );
  OAI22XL U19947 ( .A0(n16645), .A1(n32974), .B0(n32971), .B1(n26853), .Y(
        n14223) );
  OAI22XL U19948 ( .A0(n16645), .A1(n32971), .B0(n32970), .B1(n26853), .Y(
        n14224) );
  OAI22XL U19949 ( .A0(n16645), .A1(n32970), .B0(n32969), .B1(n26853), .Y(
        n14225) );
  OAI22XL U19950 ( .A0(n16645), .A1(n32969), .B0(n32968), .B1(n26853), .Y(
        n14226) );
  OAI22XL U19951 ( .A0(n16650), .A1(n32472), .B0(n32476), .B1(n26853), .Y(
        n14329) );
  OAI22XL U19952 ( .A0(n16650), .A1(n32476), .B0(n32503), .B1(n26853), .Y(
        n14330) );
  OAI22XL U19953 ( .A0(n16650), .A1(n32503), .B0(n32502), .B1(n26853), .Y(
        n14331) );
  OAI22XL U19954 ( .A0(n16650), .A1(n32502), .B0(n32501), .B1(n26853), .Y(
        n14332) );
  OAI22XL U19955 ( .A0(n16650), .A1(n32501), .B0(n32510), .B1(n26853), .Y(
        n14333) );
  OAI22XL U19956 ( .A0(n16650), .A1(n32510), .B0(n32509), .B1(n26853), .Y(
        n14334) );
  OAI22XL U19957 ( .A0(n16650), .A1(n32509), .B0(n32506), .B1(n26853), .Y(
        n14335) );
  OAI22XL U19958 ( .A0(n16650), .A1(n32506), .B0(n32514), .B1(n26853), .Y(
        n14336) );
  OAI22XL U19959 ( .A0(n16650), .A1(n32514), .B0(n32516), .B1(n26853), .Y(
        n14337) );
  OAI22XL U19960 ( .A0(n16650), .A1(n32516), .B0(n32515), .B1(n26853), .Y(
        n14338) );
  OAI22XL U19961 ( .A0(n16650), .A1(n32515), .B0(n32499), .B1(n26853), .Y(
        n14339) );
  OAI22XL U19962 ( .A0(n32491), .A1(n32499), .B0(n32490), .B1(n26853), .Y(
        n14340) );
  OAI22XL U19963 ( .A0(n32491), .A1(n32490), .B0(n32484), .B1(n26853), .Y(
        n14341) );
  OAI22XL U19964 ( .A0(n32491), .A1(n32484), .B0(n32483), .B1(n26853), .Y(
        n14342) );
  OAI22XL U19965 ( .A0(n32491), .A1(n32483), .B0(n32478), .B1(n26853), .Y(
        n14343) );
  OAI22XL U19966 ( .A0(n32491), .A1(n32478), .B0(n32473), .B1(n26853), .Y(
        n14344) );
  OAI22XL U19967 ( .A0(n32491), .A1(n32473), .B0(n32461), .B1(n26853), .Y(
        n14345) );
  OAI22XL U19968 ( .A0(n32491), .A1(n32461), .B0(n32464), .B1(n26853), .Y(
        n14346) );
  OAI22XL U19969 ( .A0(n32491), .A1(n32464), .B0(n32463), .B1(n26853), .Y(
        n14347) );
  OAI22XL U19970 ( .A0(n16650), .A1(n32749), .B0(n32748), .B1(n26853), .Y(
        n14386) );
  OAI22XL U19971 ( .A0(n16650), .A1(n32751), .B0(n32750), .B1(n26853), .Y(
        n14394) );
  OAI22XL U19972 ( .A0(n16650), .A1(n32482), .B0(n32481), .B1(n26853), .Y(
        n14451) );
  OAI22XL U19973 ( .A0(n16650), .A1(n32481), .B0(n32477), .B1(n26853), .Y(
        n14452) );
  OAI22XL U19974 ( .A0(n16650), .A1(n32477), .B0(n32467), .B1(n26853), .Y(
        n14453) );
  OAI22XL U19975 ( .A0(n16650), .A1(n32467), .B0(n32460), .B1(n26853), .Y(
        n14454) );
  OAI22XL U19976 ( .A0(n16650), .A1(n32460), .B0(n32462), .B1(n26853), .Y(
        n14455) );
  OAI22XL U19977 ( .A0(n32491), .A1(n32462), .B0(n32471), .B1(n26853), .Y(
        n14456) );
  OAI22XL U19978 ( .A0(n32491), .A1(n32471), .B0(n32487), .B1(n26853), .Y(
        n14457) );
  OAI22XL U19979 ( .A0(n32491), .A1(n32487), .B0(n32486), .B1(n26853), .Y(
        n14458) );
  OAI22XL U19980 ( .A0(n32491), .A1(n32486), .B0(n32480), .B1(n26853), .Y(
        n14459) );
  OAI22XL U19981 ( .A0(n16650), .A1(n32480), .B0(n32479), .B1(n26853), .Y(
        n14460) );
  OAI22XL U19982 ( .A0(n16650), .A1(n32479), .B0(n32496), .B1(n26853), .Y(
        n14461) );
  OAI22XL U19983 ( .A0(n16650), .A1(n32496), .B0(n32495), .B1(n26853), .Y(
        n14462) );
  OAI22XL U19984 ( .A0(n16650), .A1(n32495), .B0(n32470), .B1(n26853), .Y(
        n14463) );
  OAI22XL U19985 ( .A0(n16650), .A1(n32470), .B0(n32485), .B1(n26853), .Y(
        n14464) );
  OAI22XL U19986 ( .A0(n16650), .A1(n32485), .B0(n32489), .B1(n26853), .Y(
        n14465) );
  OAI22XL U19987 ( .A0(n16650), .A1(n32489), .B0(n32488), .B1(n26853), .Y(
        n14466) );
  OAI22XL U19988 ( .A0(n16650), .A1(n32488), .B0(n32469), .B1(n26853), .Y(
        n14467) );
  OAI22XL U19989 ( .A0(n16650), .A1(n32469), .B0(n32468), .B1(n26853), .Y(
        n14468) );
  OAI22XL U19990 ( .A0(n16650), .A1(n32466), .B0(n32465), .B1(n26853), .Y(
        n14470) );
  OAI22XL U19991 ( .A0(n16650), .A1(n32465), .B0(n32475), .B1(n26853), .Y(
        n14471) );
  OAI22XL U19992 ( .A0(n16650), .A1(n32475), .B0(n32474), .B1(n26853), .Y(
        n14472) );
  OAI22XL U19993 ( .A0(n16650), .A1(n32474), .B0(n32505), .B1(n26853), .Y(
        n14473) );
  OAI22XL U19994 ( .A0(n31084), .A1(n32505), .B0(n32508), .B1(n26853), .Y(
        n14474) );
  OAI22XL U19995 ( .A0(n16645), .A1(n32508), .B0(n32507), .B1(n26853), .Y(
        n14475) );
  OAI22XL U19996 ( .A0(n16650), .A1(n32507), .B0(n32504), .B1(n26853), .Y(
        n14476) );
  OAI22XL U19997 ( .A0(n32491), .A1(n32504), .B0(n32513), .B1(n26853), .Y(
        n14477) );
  OAI22XL U19998 ( .A0(n16650), .A1(n32513), .B0(n32512), .B1(n26853), .Y(
        n14478) );
  OAI22XL U19999 ( .A0(n31084), .A1(n32512), .B0(n32511), .B1(n26853), .Y(
        n14479) );
  OAI22XL U20000 ( .A0(n16650), .A1(n32511), .B0(n32500), .B1(n26853), .Y(
        n14480) );
  OAI22XL U20001 ( .A0(n32491), .A1(n32500), .B0(n32498), .B1(n26853), .Y(
        n14481) );
  OAI22XL U20002 ( .A0(n31077), .A1(n32498), .B0(n32497), .B1(n26853), .Y(
        n14482) );
  OAI22XL U20003 ( .A0(n16650), .A1(n32497), .B0(n32494), .B1(n26853), .Y(
        n14483) );
  OAI22XL U20004 ( .A0(n32491), .A1(n32494), .B0(n32493), .B1(n26853), .Y(
        n14484) );
  OAI22XL U20005 ( .A0(n32491), .A1(n32493), .B0(n32492), .B1(n26853), .Y(
        n14485) );
  OAI2BB2XL U20006 ( .B0(n33365), .B1(n33364), .A0N(n33365), .A1N(n33364), .Y(
        n33366) );
  XOR2XL U20007 ( .A(affine_2[15]), .B(n33362), .Y(n33365) );
  OAI2BB2XL U20008 ( .B0(n33348), .B1(n33347), .A0N(n33348), .A1N(n33347), .Y(
        n33349) );
  OAI2BB2XL U20009 ( .B0(n33338), .B1(n33337), .A0N(n33338), .A1N(n33337), .Y(
        n33339) );
  XOR2XL U20010 ( .A(affine_2[47]), .B(n33335), .Y(n33338) );
  AOI2BB2XL U20011 ( .B0(n36120), .B1(n36121), .A0N(filter_1[5]), .A1N(n36120), 
        .Y(n14664) );
  AOI2BB2XL U20012 ( .B0(n36120), .B1(n36119), .A0N(filter_1[4]), .A1N(n36120), 
        .Y(n14673) );
  AOI2BB2XL U20013 ( .B0(n36120), .B1(n36118), .A0N(filter_1[3]), .A1N(n36120), 
        .Y(n14682) );
  AOI2BB2XL U20014 ( .B0(n36120), .B1(n36117), .A0N(filter_1[2]), .A1N(n36120), 
        .Y(n14691) );
  AOI2BB2XL U20015 ( .B0(n36120), .B1(n36116), .A0N(filter_1[1]), .A1N(n36120), 
        .Y(n14700) );
  AOI2BB2XL U20016 ( .B0(n36120), .B1(n36115), .A0N(filter_1[0]), .A1N(n36120), 
        .Y(n14709) );
  AOI2BB2XL U20017 ( .B0(n34813), .B1(n34812), .A0N(pool[21]), .A1N(n34813), 
        .Y(N29237) );
  AOI2BB2XL U20018 ( .B0(n34841), .B1(n34840), .A0N(n34840), .A1N(pool[36]), 
        .Y(N29252) );
  AOI2BB2XL U20019 ( .B0(n34791), .B1(n34790), .A0N(pool[1]), .A1N(n34791), 
        .Y(N29217) );
  AOI2BB2XL U20020 ( .B0(n34818), .B1(n34817), .A0N(n34817), .A1N(pool[26]), 
        .Y(N29242) );
  AOI2BB2XL U20021 ( .B0(n34803), .B1(n34802), .A0N(n34802), .A1N(pool[11]), 
        .Y(N29227) );
  AOI2BB2XL U20022 ( .B0(n34857), .B1(n34861), .A0N(n34861), .A1N(pool[41]), 
        .Y(N29257) );
  AOI2BB2XL U20023 ( .B0(n34836), .B1(n34835), .A0N(n34835), .A1N(pool[31]), 
        .Y(N29247) );
  NOR2XL U20024 ( .A(n23820), .B(n16655), .Y(n23821) );
  AOI2BB2XL U20025 ( .B0(n36114), .B1(n36113), .A0N(filter_1_bias[1]), .A1N(
        n36114), .Y(n14718) );
  AOI2BB2XL U20026 ( .B0(n34888), .B1(n34887), .A0N(pool[66]), .A1N(n34888), 
        .Y(N29282) );
  AOI2BB2XL U20027 ( .B0(n34868), .B1(n34872), .A0N(n34872), .A1N(pool[51]), 
        .Y(N29267) );
  AOI2BB2XL U20028 ( .B0(n34893), .B1(n34892), .A0N(n34892), .A1N(pool[71]), 
        .Y(N29287) );
  AOI2BB2XL U20029 ( .B0(n34875), .B1(n34874), .A0N(n34874), .A1N(pool[56]), 
        .Y(N29272) );
  AOI2BB2XL U20030 ( .B0(n34898), .B1(n34897), .A0N(n34897), .A1N(pool[76]), 
        .Y(N29292) );
  AOI2BB1XL U20031 ( .A0N(n34237), .A1N(n36091), .B0(n34236), .Y(n34238) );
  NOR2X1 U20032 ( .A(n34237), .B(n34235), .Y(n34234) );
  NOR2X1 U20033 ( .A(n29770), .B(n29769), .Y(n29772) );
  AOI2BB2XL U20034 ( .B0(n35011), .B1(n35015), .A0N(n35015), .A1N(pool[111]), 
        .Y(N29327) );
  AOI2BB2XL U20035 ( .B0(n35023), .B1(n35027), .A0N(n35027), .A1N(pool[126]), 
        .Y(N29342) );
  AOI2BB2XL U20036 ( .B0(n34975), .B1(n34979), .A0N(n34979), .A1N(pool[96]), 
        .Y(N29312) );
  AOI2BB2XL U20037 ( .B0(n35017), .B1(n35018), .A0N(n35018), .A1N(pool[116]), 
        .Y(N29332) );
  AOI2BB2XL U20038 ( .B0(n35001), .B1(n34996), .A0N(n34995), .A1N(n35001), .Y(
        N29317) );
  AOI2BB2XL U20039 ( .B0(n35010), .B1(n35005), .A0N(n35004), .A1N(n35010), .Y(
        N29322) );
  AOI2BB2XL U20040 ( .B0(n35247), .B1(n35252), .A0N(n35252), .A1N(pool[131]), 
        .Y(N29347) );
  NOR2X1 U20041 ( .A(n30525), .B(n30524), .Y(n30527) );
  NOR2X1 U20042 ( .A(n30538), .B(n30537), .Y(n30540) );
  AOI2BB2XL U20043 ( .B0(n34816), .B1(n34815), .A0N(n34815), .A1N(n34814), .Y(
        N29238) );
  AOI2BB2XL U20044 ( .B0(n34844), .B1(n34843), .A0N(n34842), .A1N(n34844), .Y(
        N29253) );
  AOI2BB2XL U20045 ( .B0(n34801), .B1(n34800), .A0N(n34800), .A1N(n34799), .Y(
        N29223) );
  AOI2BB2XL U20046 ( .B0(n34793), .B1(n34795), .A0N(n34795), .A1N(n34792), .Y(
        N29218) );
  AOI2BB2XL U20047 ( .B0(n34811), .B1(n34810), .A0N(n34810), .A1N(n34809), .Y(
        N29233) );
  AOI2BB2XL U20048 ( .B0(n34860), .B1(n34859), .A0N(n34858), .A1N(n34860), .Y(
        N29258) );
  AOI2BB2XL U20049 ( .B0(n34839), .B1(n34838), .A0N(n34837), .A1N(n34839), .Y(
        N29248) );
  NOR2X1 U20050 ( .A(n30461), .B(n30460), .Y(n30463) );
  NOR2X1 U20051 ( .A(n27374), .B(n27373), .Y(n27376) );
  AOI31XL U20052 ( .A0(n36056), .A1(n33541), .A2(n33540), .B0(conv_1[422]), 
        .Y(n33543) );
  AOI2BB2XL U20053 ( .B0(n36114), .B1(n36112), .A0N(filter_1_bias[2]), .A1N(
        n36114), .Y(n14721) );
  AOI2BB2XL U20054 ( .B0(n34891), .B1(n34890), .A0N(n34890), .A1N(n34889), .Y(
        N29283) );
  AOI2BB2XL U20055 ( .B0(n34871), .B1(n34870), .A0N(n34869), .A1N(n34871), .Y(
        N29268) );
  AOI2BB2XL U20056 ( .B0(n34867), .B1(n34866), .A0N(n34866), .A1N(n34865), .Y(
        N29263) );
  AOI2BB2XL U20057 ( .B0(n34880), .B1(n34877), .A0N(n34876), .A1N(n34880), .Y(
        N29273) );
  AOI2BB2XL U20058 ( .B0(n34941), .B1(n34940), .A0N(n34940), .A1N(n34939), .Y(
        N29303) );
  AOI2BB1XL U20059 ( .A0N(n34620), .A1N(n35902), .B0(n34619), .Y(n34622) );
  NOR2X1 U20060 ( .A(n34620), .B(n34618), .Y(n34617) );
  AOI2BB2XL U20061 ( .B0(n35014), .B1(n35013), .A0N(n35012), .A1N(n35014), .Y(
        N29328) );
  AOI2BB2XL U20062 ( .B0(n35026), .B1(n35025), .A0N(n35024), .A1N(n35026), .Y(
        N29343) );
  AOI2BB2XL U20063 ( .B0(n34978), .B1(n34977), .A0N(n34976), .A1N(n34978), .Y(
        N29313) );
  AOI2BB2XL U20064 ( .B0(n34946), .B1(n34945), .A0N(n34945), .A1N(n34944), .Y(
        N29308) );
  AOI2BB2XL U20065 ( .B0(n34998), .B1(n34997), .A0N(n34997), .A1N(pool[102]), 
        .Y(N29318) );
  AOI2BB2XL U20066 ( .B0(n35007), .B1(n35006), .A0N(n35006), .A1N(pool[107]), 
        .Y(N29323) );
  AOI2BB2XL U20067 ( .B0(n35250), .B1(n35249), .A0N(n35248), .A1N(n35250), .Y(
        N29348) );
  NOR2X1 U20068 ( .A(n30513), .B(n30512), .Y(n30515) );
  AOI2BB1XL U20069 ( .A0N(n34611), .A1N(n35610), .B0(n34610), .Y(n34612) );
  NOR2X1 U20070 ( .A(n34611), .B(n34609), .Y(n34608) );
  NOR2X1 U20071 ( .A(n30551), .B(n30550), .Y(n30553) );
  AOI2BB2XL U20072 ( .B0(n34862), .B1(n34861), .A0N(n34861), .A1N(pool[43]), 
        .Y(N29259) );
  NOR2X1 U20073 ( .A(n24688), .B(n24690), .Y(n23470) );
  AOI2BB2XL U20074 ( .B0(n36114), .B1(n36111), .A0N(filter_1_bias[3]), .A1N(
        n36114), .Y(n14724) );
  AOI2BB2XL U20075 ( .B0(n34873), .B1(n34872), .A0N(n34872), .A1N(pool[53]), 
        .Y(N29269) );
  AOI2BB2XL U20076 ( .B0(n34943), .B1(n34942), .A0N(pool[88]), .A1N(n34943), 
        .Y(N29304) );
  AOI2BB1XL U20077 ( .A0N(n34104), .A1N(n36091), .B0(n34103), .Y(n34106) );
  NOR2X1 U20078 ( .A(n34104), .B(n34102), .Y(n34101) );
  NOR2X1 U20079 ( .A(n29554), .B(n29553), .Y(n29556) );
  NOR2X1 U20080 ( .A(n27701), .B(n27703), .Y(n23797) );
  NOR2X1 U20081 ( .A(n27551), .B(n27552), .Y(n23583) );
  AOI2BB2XL U20082 ( .B0(n35016), .B1(n35015), .A0N(n35015), .A1N(pool[113]), 
        .Y(N29329) );
  AOI2BB2XL U20083 ( .B0(n35028), .B1(n35027), .A0N(n35027), .A1N(pool[128]), 
        .Y(N29344) );
  AOI2BB2XL U20084 ( .B0(n34980), .B1(n34979), .A0N(n34979), .A1N(pool[98]), 
        .Y(N29314) );
  AOI2BB2XL U20085 ( .B0(n34948), .B1(n34947), .A0N(pool[93]), .A1N(n34948), 
        .Y(N29309) );
  AOI2BB2XL U20086 ( .B0(n35019), .B1(n35018), .A0N(n35018), .A1N(pool[118]), 
        .Y(N29334) );
  AOI2BB2XL U20087 ( .B0(n35001), .B1(n35000), .A0N(n34999), .A1N(n35001), .Y(
        N29319) );
  AOI2BB2XL U20088 ( .B0(n35010), .B1(n35009), .A0N(n35008), .A1N(n35010), .Y(
        N29324) );
  AOI2BB2XL U20089 ( .B0(n35251), .B1(n35252), .A0N(n35252), .A1N(pool[133]), 
        .Y(N29349) );
  NOR2X1 U20090 ( .A(n30185), .B(n30184), .Y(n30187) );
  NOR2X1 U20091 ( .A(n29415), .B(n29414), .Y(n29417) );
  NOR2X1 U20092 ( .A(n29670), .B(n29669), .Y(n29672) );
  AOI2BB1XL U20093 ( .A0N(n34112), .A1N(n35598), .B0(n34111), .Y(n34113) );
  NOR2X1 U20094 ( .A(n34112), .B(n34110), .Y(n34109) );
  AOI2BB2XL U20095 ( .B0(n34796), .B1(n34795), .A0N(n34795), .A1N(n34794), .Y(
        N29220) );
  NOR2X1 U20096 ( .A(n30696), .B(n30695), .Y(n30698) );
  NOR2X1 U20097 ( .A(n27399), .B(n27398), .Y(n27401) );
  NOR2X1 U20098 ( .A(n27007), .B(n27006), .Y(n27009) );
  NOR2X1 U20099 ( .A(n27393), .B(n27392), .Y(n27395) );
  NOR2X1 U20100 ( .A(n23910), .B(n23909), .Y(n23912) );
  AOI2BB2XL U20101 ( .B0(n36114), .B1(n36110), .A0N(filter_1_bias[4]), .A1N(
        n36114), .Y(n14727) );
  AOI2BB2XL U20102 ( .B0(n34880), .B1(n34879), .A0N(n34878), .A1N(n34880), .Y(
        N29275) );
  NOR2X1 U20103 ( .A(n29029), .B(n29028), .Y(n29031) );
  NOR2X1 U20104 ( .A(n29017), .B(n29016), .Y(n29019) );
  NOR2X1 U20105 ( .A(n28877), .B(n28876), .Y(n28879) );
  AOI2BB1XL U20106 ( .A0N(n34407), .A1N(n35894), .B0(n34406), .Y(n34409) );
  NOR2X1 U20107 ( .A(n25280), .B(n25278), .Y(n25277) );
  NOR2X1 U20108 ( .A(n29714), .B(n29713), .Y(n29716) );
  AOI2BB2XL U20109 ( .B0(n35253), .B1(n35252), .A0N(n35252), .A1N(pool[134]), 
        .Y(N29350) );
  AOI32XL U20110 ( .A0(n36056), .A1(n34096), .A2(n34095), .B0(conv_3[499]), 
        .B1(n34094), .Y(n34098) );
  NOR2X1 U20111 ( .A(n22191), .B(n22190), .Y(n22193) );
  AOI32XL U20112 ( .A0(n36056), .A1(n34076), .A2(n34075), .B0(conv_3[424]), 
        .B1(n34074), .Y(n34077) );
  NOR2X1 U20113 ( .A(n31404), .B(n31405), .Y(n23225) );
  NOR2X1 U20114 ( .A(n26152), .B(n26153), .Y(n22166) );
  NOR2X1 U20115 ( .A(n26524), .B(n26525), .Y(n23625) );
  NOR2X1 U20116 ( .A(n31666), .B(n31667), .Y(n22879) );
  NOR2X1 U20117 ( .A(n23700), .B(n23698), .Y(n23697) );
  AOI211XL U20118 ( .A0(n34963), .A1(n28406), .B0(n25311), .C0(n25310), .Y(
        n25436) );
  NOR2X1 U20119 ( .A(n34833), .B(n34832), .Y(n34834) );
  NOR2X1 U20120 ( .A(n24917), .B(n24915), .Y(n24914) );
  NOR2X1 U20121 ( .A(n26339), .B(n26337), .Y(n26336) );
  NOR2X1 U20122 ( .A(n30324), .B(n33209), .Y(n29975) );
  AOI2BB1XL U20123 ( .A0N(n29828), .A1N(n33506), .B0(n29827), .Y(n29829) );
  NOR2X1 U20124 ( .A(n29828), .B(n29826), .Y(n29825) );
  NOR2X1 U20125 ( .A(n26346), .B(n26344), .Y(n26343) );
  NOR2X1 U20126 ( .A(n27244), .B(n27243), .Y(n27246) );
  NOR2X1 U20127 ( .A(n25236), .B(n25234), .Y(n25233) );
  AOI31XL U20128 ( .A0(n36056), .A1(n27582), .A2(n27581), .B0(n35549), .Y(
        n27587) );
  OAI21XL U20129 ( .A0(n34776), .A1(n34775), .B0(n34774), .Y(n34777) );
  NOR2X1 U20130 ( .A(n29299), .B(n29298), .Y(n29301) );
  NOR2X1 U20131 ( .A(n26520), .B(n25255), .Y(n25254) );
  AOI31XL U20132 ( .A0(n36056), .A1(n35480), .A2(n35479), .B0(n35549), .Y(
        n35481) );
  NOR2X1 U20133 ( .A(n33654), .B(n33653), .Y(n33650) );
  NOR2X1 U20134 ( .A(n29275), .B(n29274), .Y(n29277) );
  NOR2X1 U20135 ( .A(n34340), .B(n34338), .Y(n34337) );
  AOI2BB1XL U20136 ( .A0N(n34311), .A1N(n35458), .B0(n34310), .Y(n34312) );
  NOR2X1 U20137 ( .A(n34311), .B(n34309), .Y(n34308) );
  AOI2BB1XL U20138 ( .A0N(n34287), .A1N(n35458), .B0(n34286), .Y(n34288) );
  NOR2X1 U20139 ( .A(n34287), .B(n34285), .Y(n34284) );
  AOI2BB1XL U20140 ( .A0N(n35455), .A1N(n31362), .B0(n31364), .Y(n23153) );
  AOI32XL U20141 ( .A0(n35458), .A1(n27580), .A2(n27579), .B0(n27578), .B1(
        n27580), .Y(n16096) );
  AOI31XL U20142 ( .A0(n36056), .A1(n27575), .A2(n27574), .B0(n35549), .Y(
        n27580) );
  NAND2XL U20143 ( .A(conv_1[374]), .B(n33132), .Y(n33131) );
  NOR2X1 U20144 ( .A(n33889), .B(n33887), .Y(n33886) );
  AOI2BB1XL U20145 ( .A0N(n34255), .A1N(n34263), .B0(n34254), .Y(n34256) );
  NOR2X1 U20146 ( .A(n34255), .B(n34253), .Y(n34252) );
  AOI2BB1XL U20147 ( .A0N(n34264), .A1N(n34263), .B0(n34262), .Y(n34265) );
  NOR2X1 U20148 ( .A(n34264), .B(n34261), .Y(n34260) );
  NOR2X1 U20149 ( .A(n23310), .B(n23309), .Y(n23312) );
  NOR2X1 U20150 ( .A(n25287), .B(n25285), .Y(n25284) );
  AOI2BB1XL U20151 ( .A0N(n34326), .A1N(n34325), .B0(n34324), .Y(n34327) );
  NOR2X1 U20152 ( .A(n34326), .B(n34323), .Y(n34322) );
  AOI2BB1XL U20153 ( .A0N(n34317), .A1N(n34325), .B0(n34316), .Y(n34318) );
  NOR2X1 U20154 ( .A(n34317), .B(n34315), .Y(n34314) );
  NOR2X1 U20155 ( .A(n29311), .B(n29310), .Y(n29313) );
  AOI31XL U20156 ( .A0(n36056), .A1(n35429), .A2(n35428), .B0(n35549), .Y(
        n35430) );
  AOI32XL U20157 ( .A0(n36056), .A1(n34083), .A2(n34082), .B0(conv_1[268]), 
        .B1(n34081), .Y(n34084) );
  AOI31XL U20158 ( .A0(n36056), .A1(n29197), .A2(n27563), .B0(n35549), .Y(
        n27566) );
  AOI32XL U20159 ( .A0(n36056), .A1(n27561), .A2(n24695), .B0(conv_1[260]), 
        .B1(n24694), .Y(n24696) );
  NOR2X1 U20160 ( .A(n27562), .B(n27560), .Y(n24695) );
  AOI32XL U20161 ( .A0(n36056), .A1(n27981), .A2(n26974), .B0(conv_1[253]), 
        .B1(n26973), .Y(n26975) );
  NOR2X1 U20162 ( .A(n33663), .B(n33662), .Y(n33659) );
  NOR2X1 U20163 ( .A(n26970), .B(n26971), .Y(n26495) );
  AOI2BB1XL U20164 ( .A0N(n34333), .A1N(n35417), .B0(n34332), .Y(n34334) );
  NOR2X1 U20165 ( .A(n34333), .B(n34331), .Y(n34330) );
  AOI2BB1XL U20166 ( .A0N(n34280), .A1N(n35408), .B0(n34279), .Y(n34282) );
  AOI2BB1XL U20167 ( .A0N(n34304), .A1N(n35395), .B0(n34303), .Y(n34305) );
  AOI32XL U20168 ( .A0(n36056), .A1(n25441), .A2(n25440), .B0(conv_1[221]), 
        .B1(n25439), .Y(n25442) );
  NOR2X1 U20169 ( .A(n34543), .B(n34541), .Y(n34540) );
  NOR2X1 U20170 ( .A(n24684), .B(n24682), .Y(n24681) );
  AOI2BB1XL U20171 ( .A0N(n34064), .A1N(n35384), .B0(n34063), .Y(n34065) );
  NOR2X1 U20172 ( .A(n34064), .B(n34062), .Y(n34061) );
  NOR2X1 U20173 ( .A(n35379), .B(n23682), .Y(n23679) );
  NOR2X1 U20174 ( .A(n23445), .B(n23444), .Y(n23441) );
  AOI32XL U20175 ( .A0(n36056), .A1(n34122), .A2(n34121), .B0(conv_1[193]), 
        .B1(n34120), .Y(n34123) );
  NAND2XL U20176 ( .A(n34119), .B(n34118), .Y(n34121) );
  AOI2BB1XL U20177 ( .A0N(n34090), .A1N(n35368), .B0(n34089), .Y(n34091) );
  NOR2X1 U20178 ( .A(n34090), .B(n34088), .Y(n34087) );
  AOI2BB1XL U20179 ( .A0N(n35365), .A1N(n35364), .B0(n35363), .Y(n35366) );
  AOI2BB1XL U20180 ( .A0N(n34049), .A1N(n34048), .B0(n34047), .Y(n34050) );
  NOR2X1 U20181 ( .A(n34049), .B(n34046), .Y(n34045) );
  NOR2X1 U20182 ( .A(n23400), .B(n23399), .Y(n23402) );
  AOI2BB1XL U20183 ( .A0N(n34272), .A1N(n34271), .B0(n34270), .Y(n34273) );
  NOR2X1 U20184 ( .A(n34272), .B(n34269), .Y(n34268) );
  NOR2X1 U20185 ( .A(n25452), .B(n25450), .Y(n25449) );
  AOI2BB1XL U20186 ( .A0N(n34297), .A1N(n34296), .B0(n34295), .Y(n34298) );
  OAI2BB1XL U20187 ( .A0N(n33912), .A1N(n33491), .B0(n34296), .Y(n33492) );
  AOI32XL U20188 ( .A0(n36056), .A1(n33242), .A2(n33241), .B0(conv_1[118]), 
        .B1(n33240), .Y(n33243) );
  NAND2XL U20189 ( .A(n33239), .B(n33238), .Y(n33241) );
  NOR2X1 U20190 ( .A(n25096), .B(n25094), .Y(n25093) );
  NOR2X1 U20191 ( .A(n29293), .B(n29292), .Y(n29295) );
  AOI2BB1XL U20192 ( .A0N(n31336), .A1N(n31361), .B0(n26844), .Y(n26845) );
  NOR2X1 U20193 ( .A(n31336), .B(n26843), .Y(n26842) );
  AOI32XL U20194 ( .A0(n36056), .A1(n26777), .A2(n26517), .B0(conv_1[95]), 
        .B1(n26516), .Y(n26518) );
  OAI211XL U20195 ( .A0(n34676), .A1(n31341), .B0(n16652), .C0(n31340), .Y(
        n16359) );
  NOR2X1 U20196 ( .A(n26736), .B(n24928), .Y(n24927) );
  AOI2BB1XL U20197 ( .A0N(n34058), .A1N(n34057), .B0(n34056), .Y(n34059) );
  NOR2X1 U20198 ( .A(n34058), .B(n34055), .Y(n34054) );
  NOR2X1 U20199 ( .A(n24936), .B(n24934), .Y(n24933) );
  AOI2BB1XL U20200 ( .A0N(n26310), .A1N(n35327), .B0(n26144), .Y(n26145) );
  NOR2X1 U20201 ( .A(n26310), .B(n26143), .Y(n26142) );
  NOR2X1 U20202 ( .A(n33638), .B(n33637), .Y(n33634) );
  NOR2X1 U20203 ( .A(n33638), .B(n27201), .Y(n27198) );
  AOI31XL U20204 ( .A0(n36056), .A1(n32518), .A2(n32519), .B0(n35549), .Y(
        n32524) );
  OR2XL U20205 ( .A(n35549), .B(n35313), .Y(n16409) );
  OAI21XL U20206 ( .A0(n33251), .A1(n35289), .B0(n33250), .Y(n33252) );
  OAI2BB1XL U20207 ( .A0N(conv_1[41]), .A1N(n35306), .B0(n35305), .Y(n16422)
         );
  AOI31XL U20208 ( .A0(n36056), .A1(n35304), .A2(n35303), .B0(n35549), .Y(
        n35305) );
  AOI32XL U20209 ( .A0(n36056), .A1(n27333), .A2(n26507), .B0(conv_1[20]), 
        .B1(n26506), .Y(n26508) );
  AOI32XL U20210 ( .A0(n36056), .A1(n27362), .A2(n26300), .B0(conv_1[13]), 
        .B1(n26299), .Y(n26301) );
  NOR2X1 U20211 ( .A(n34553), .B(n34550), .Y(n34549) );
  AOI2BB2XL U20212 ( .B0(n36114), .B1(n36109), .A0N(filter_1_bias[5]), .A1N(
        n36114), .Y(n14730) );
  NOR2X1 U20213 ( .A(n33629), .B(n33373), .Y(n33370) );
  NOR2X1 U20214 ( .A(n29629), .B(n29627), .Y(n29626) );
  MXI2XL U20215 ( .A(n34923), .B(n34922), .S0(n34926), .Y(N29296) );
  AOI2BB1XL U20216 ( .A0N(n31014), .A1N(n31013), .B0(n31012), .Y(n31015) );
  NOR2X1 U20217 ( .A(n31014), .B(n31011), .Y(n31010) );
  AOI2BB1XL U20218 ( .A0N(n33580), .A1N(n27794), .B0(n27793), .Y(n27796) );
  NOR2X1 U20219 ( .A(n27776), .B(n27775), .Y(n27778) );
  OAI211XL U20220 ( .A0(n34520), .A1(n29443), .B0(n34669), .C0(n29442), .Y(
        n14854) );
  NAND2XL U20221 ( .A(conv_2[524]), .B(n29441), .Y(n29440) );
  AOI22XL U20222 ( .A0(conv_2[523]), .A1(n29439), .B0(n29438), .B1(n29437), 
        .Y(n29441) );
  NOR2X1 U20223 ( .A(n33168), .B(n30913), .Y(n30912) );
  OR2XL U20224 ( .A(n16651), .B(n36078), .Y(n14870) );
  AOI2BB1XL U20225 ( .A0N(n34178), .A1N(n34177), .B0(n34176), .Y(n34179) );
  NOR2X1 U20226 ( .A(n34178), .B(n34175), .Y(n34174) );
  NOR2X1 U20227 ( .A(n27872), .B(n27873), .Y(n27869) );
  AOI2BB1XL U20228 ( .A0N(n33896), .A1N(n34177), .B0(n33895), .Y(n33897) );
  NOR2X1 U20229 ( .A(n33896), .B(n33894), .Y(n33893) );
  NOR2X1 U20230 ( .A(n30881), .B(n30879), .Y(n30878) );
  AOI32XL U20231 ( .A0(n36056), .A1(n34734), .A2(n34733), .B0(conv_2[448]), 
        .B1(n34732), .Y(n34736) );
  NOR2X1 U20232 ( .A(n30966), .B(n30964), .Y(n30963) );
  NOR2X1 U20233 ( .A(n30870), .B(n30868), .Y(n30867) );
  OR2XL U20234 ( .A(n16651), .B(n36064), .Y(n14912) );
  AOI2BB1XL U20235 ( .A0N(n34207), .A1N(n36053), .B0(n34206), .Y(n34208) );
  AOI2BB1XL U20236 ( .A0N(n34215), .A1N(n36053), .B0(n34214), .Y(n34216) );
  NOR2X1 U20237 ( .A(n34215), .B(n34213), .Y(n34212) );
  AOI32XL U20238 ( .A0(n36056), .A1(n34040), .A2(n34039), .B0(conv_2[418]), 
        .B1(n34038), .Y(n34041) );
  NAND2XL U20239 ( .A(n34037), .B(n34036), .Y(n34039) );
  AOI31XL U20240 ( .A0(n36056), .A1(n36049), .A2(n36048), .B0(n16651), .Y(
        n36050) );
  NOR2X1 U20241 ( .A(n36038), .B(n36037), .Y(n36039) );
  NOR2X1 U20242 ( .A(n36045), .B(n33691), .Y(n33688) );
  NOR2X1 U20243 ( .A(n34640), .B(n34638), .Y(n34637) );
  NOR2X1 U20244 ( .A(n28115), .B(n28114), .Y(n28117) );
  NOR2X1 U20245 ( .A(n28013), .B(n28012), .Y(n28015) );
  NOR2X1 U20246 ( .A(n29445), .B(n29444), .Y(n29447) );
  AOI2BB1XL U20247 ( .A0N(n34576), .A1N(n36017), .B0(n34575), .Y(n34577) );
  AOI2BB1XL U20248 ( .A0N(n34568), .A1N(n36017), .B0(n34567), .Y(n34569) );
  NOR2X1 U20249 ( .A(n34568), .B(n34566), .Y(n34565) );
  NOR2X1 U20250 ( .A(n33931), .B(n33929), .Y(n33928) );
  NOR2X1 U20251 ( .A(n29615), .B(n29613), .Y(n29612) );
  AOI2BB1XL U20252 ( .A0N(n33938), .A1N(n35986), .B0(n33937), .Y(n33939) );
  NOR2X1 U20253 ( .A(n28058), .B(n26354), .Y(n26353) );
  AOI222XL U20254 ( .A0(conv_2[313]), .A1(n34025), .B0(conv_2[313]), .B1(
        n34024), .C0(n34023), .C1(n34022), .Y(n34027) );
  AOI32XL U20255 ( .A0(n36056), .A1(n30861), .A2(n30860), .B0(conv_2[305]), 
        .B1(n30859), .Y(n30862) );
  NOR2X1 U20256 ( .A(n32981), .B(n32979), .Y(n32978) );
  AOI32XL U20257 ( .A0(n36056), .A1(n30892), .A2(n30891), .B0(conv_2[290]), 
        .B1(n30890), .Y(n30893) );
  OAI211XL U20258 ( .A0(n34520), .A1(n33300), .B0(n34669), .C0(n33299), .Y(
        n15004) );
  AOI22XL U20259 ( .A0(conv_2[298]), .A1(n33296), .B0(n33295), .B1(n33294), 
        .Y(n33298) );
  AOI32XL U20260 ( .A0(n36056), .A1(n30997), .A2(n30996), .B0(conv_2[283]), 
        .B1(n30995), .Y(n30998) );
  NOR2X1 U20261 ( .A(n30990), .B(n30988), .Y(n30987) );
  NOR2X1 U20262 ( .A(n28007), .B(n28006), .Y(n28009) );
  NOR2X1 U20263 ( .A(n34600), .B(n34599), .Y(n34603) );
  NOR2X1 U20264 ( .A(n28178), .B(n28177), .Y(n28180) );
  AOI32XL U20265 ( .A0(n36056), .A1(n34148), .A2(n34147), .B0(conv_2[253]), 
        .B1(n34146), .Y(n34149) );
  NOR2X1 U20266 ( .A(n35942), .B(n33683), .Y(n33680) );
  NOR2X1 U20267 ( .A(n30936), .B(n30934), .Y(n30933) );
  NOR2X1 U20268 ( .A(n29513), .B(n29512), .Y(n29515) );
  AOI31XL U20269 ( .A0(n36056), .A1(n30430), .A2(n28666), .B0(n16651), .Y(
        n28669) );
  AOI2BB1XL U20270 ( .A0N(n30952), .A1N(n35917), .B0(n30951), .Y(n30953) );
  NOR2X1 U20271 ( .A(n35914), .B(n33457), .Y(n33454) );
  AOI31XL U20272 ( .A0(n36056), .A1(n29891), .A2(n28656), .B0(n16651), .Y(
        n28659) );
  AOI2BB1XL U20273 ( .A0N(n34590), .A1N(n34589), .B0(n34588), .Y(n34591) );
  NOR2X1 U20274 ( .A(n34590), .B(n34587), .Y(n34586) );
  NOR2X1 U20275 ( .A(n29839), .B(n29840), .Y(n29836) );
  OAI211XL U20276 ( .A0(n33442), .A1(n34598), .B0(n34735), .C0(n34597), .Y(
        n15084) );
  NAND2XL U20277 ( .A(conv_2[179]), .B(n34596), .Y(n34595) );
  AOI32XL U20278 ( .A0(n36056), .A1(n26361), .A2(n26360), .B0(conv_2[163]), 
        .B1(n26359), .Y(n26362) );
  NAND2XL U20279 ( .A(n26358), .B(n26357), .Y(n26360) );
  AOI2BB1XL U20280 ( .A0N(n33951), .A1N(n34631), .B0(n33950), .Y(n33952) );
  NOR2X1 U20281 ( .A(n33951), .B(n33949), .Y(n33948) );
  AOI2BB1XL U20282 ( .A0N(n33944), .A1N(n34631), .B0(n33943), .Y(n33945) );
  NOR2X1 U20283 ( .A(n33944), .B(n33942), .Y(n33941) );
  AOI2BB1XL U20284 ( .A0N(n34632), .A1N(n34631), .B0(n34630), .Y(n34633) );
  NOR2X1 U20285 ( .A(n34632), .B(n34629), .Y(n34628) );
  AOI2BB1XL U20286 ( .A0N(n34362), .A1N(n35902), .B0(n34361), .Y(n34363) );
  NOR2X1 U20287 ( .A(n34362), .B(n34360), .Y(n34359) );
  AOI2BB1XL U20288 ( .A0N(n34355), .A1N(n34491), .B0(n34354), .Y(n34356) );
  NOR2X1 U20289 ( .A(n34355), .B(n34353), .Y(n34352) );
  AOI2BB1XL U20290 ( .A0N(n34348), .A1N(n34491), .B0(n34347), .Y(n34349) );
  NOR2X1 U20291 ( .A(n30062), .B(n30061), .Y(n30064) );
  NOR2X1 U20292 ( .A(n34125), .B(n34124), .Y(n34127) );
  AOI2BB1XL U20293 ( .A0N(n34368), .A1N(n35894), .B0(n34367), .Y(n34369) );
  NOR2X1 U20294 ( .A(n34368), .B(n34366), .Y(n34365) );
  NOR2X1 U20295 ( .A(n34647), .B(n34645), .Y(n34644) );
  AOI31XL U20296 ( .A0(n36056), .A1(n30137), .A2(n28681), .B0(n16651), .Y(
        n28684) );
  NOR2X1 U20297 ( .A(n28679), .B(n25681), .Y(n25680) );
  AOI32XL U20298 ( .A0(n36056), .A1(n33292), .A2(n33291), .B0(conv_2[103]), 
        .B1(n33290), .Y(n33293) );
  NOR2X1 U20299 ( .A(n30944), .B(n30942), .Y(n30941) );
  AOI32XL U20300 ( .A0(n36056), .A1(n32671), .A2(n30929), .B0(conv_2[88]), 
        .B1(n30928), .Y(n30930) );
  NAND2XL U20301 ( .A(n32673), .B(n32672), .Y(n30929) );
  NOR2X1 U20302 ( .A(n35876), .B(n33813), .Y(n33810) );
  AOI32XL U20303 ( .A0(n35879), .A1(n28746), .A2(n28745), .B0(n30174), .B1(
        n28746), .Y(n15149) );
  NOR2X1 U20304 ( .A(n30977), .B(n30975), .Y(n30974) );
  NOR2X1 U20305 ( .A(n30118), .B(n30119), .Y(n30109) );
  NOR2X1 U20306 ( .A(n33735), .B(n30107), .Y(n18975) );
  NOR2X1 U20307 ( .A(n27820), .B(n27819), .Y(n27822) );
  NOR2X1 U20308 ( .A(n27807), .B(n27806), .Y(n27804) );
  NOR2X1 U20309 ( .A(n29622), .B(n29620), .Y(n29619) );
  NOR2X1 U20310 ( .A(n33588), .B(n33587), .Y(n33584) );
  NOR2X1 U20311 ( .A(n33620), .B(n27917), .Y(n27914) );
  AOI31XL U20312 ( .A0(n36056), .A1(n28671), .A2(n28670), .B0(n16651), .Y(
        n28677) );
  NOR2X1 U20313 ( .A(n33620), .B(n33619), .Y(n33616) );
  AOI32XL U20314 ( .A0(n30412), .A1(n27559), .A2(n27558), .B0(n27832), .B1(
        n27559), .Y(n15191) );
  AOI31XL U20315 ( .A0(n36056), .A1(n27830), .A2(n27556), .B0(n16651), .Y(
        n27559) );
  NOR2X1 U20316 ( .A(n29594), .B(n29592), .Y(n29591) );
  NOR2X1 U20317 ( .A(n29587), .B(n29585), .Y(n29584) );
  AOI32XL U20318 ( .A0(n31191), .A1(n28963), .A2(n28962), .B0(n28961), .B1(
        n28963), .Y(n15389) );
  AOI32XL U20319 ( .A0(n31191), .A1(n27573), .A2(n27572), .B0(n27571), .B1(
        n27573), .Y(n15391) );
  AOI31XL U20320 ( .A0(n36056), .A1(n27568), .A2(n27567), .B0(n16653), .Y(
        n27573) );
  MXI2XL U20321 ( .A(n34974), .B(n34973), .S0(n34978), .Y(N29311) );
  MXI2XL U20322 ( .A(n34994), .B(n34993), .S0(n35001), .Y(N29316) );
  AOI32XL U20323 ( .A0(n36056), .A1(n33306), .A2(n33305), .B0(conv_3[523]), 
        .B1(n33304), .Y(n33307) );
  NOR2X1 U20324 ( .A(n26682), .B(n26680), .Y(n26679) );
  NOR2X1 U20325 ( .A(n32071), .B(n32070), .Y(n32073) );
  NOR2X1 U20326 ( .A(n33964), .B(n33962), .Y(n33961) );
  NOR2BXL U20327 ( .AN(n32340), .B(n32339), .Y(n32342) );
  NOR2X1 U20328 ( .A(n32334), .B(n32333), .Y(n32336) );
  AOI32XL U20329 ( .A0(n36056), .A1(n26124), .A2(n26123), .B0(conv_3[470]), 
        .B1(n26122), .Y(n26125) );
  NOR2X1 U20330 ( .A(n26121), .B(n26120), .Y(n26123) );
  NOR2BXL U20331 ( .AN(n31524), .B(n31523), .Y(n31526) );
  NOR2X1 U20332 ( .A(n35802), .B(n35801), .Y(n35803) );
  NOR2X1 U20333 ( .A(n33780), .B(n33779), .Y(n33775) );
  NOR2X1 U20334 ( .A(n33761), .B(n33760), .Y(n33757) );
  NOR2X1 U20335 ( .A(n33761), .B(n32110), .Y(n32107) );
  NOR2X1 U20336 ( .A(n32586), .B(n32584), .Y(n32583) );
  NOR2BXL U20337 ( .AN(n32582), .B(n32157), .Y(n31728) );
  AOI32XL U20338 ( .A0(n36056), .A1(n32579), .A2(n32578), .B0(conv_3[425]), 
        .B1(n32577), .Y(n32580) );
  NOR2X1 U20339 ( .A(n32576), .B(n32575), .Y(n32578) );
  NOR2X1 U20340 ( .A(n32011), .B(n32010), .Y(n32013) );
  NOR2X1 U20341 ( .A(n32563), .B(n32561), .Y(n32560) );
  AOI32XL U20342 ( .A0(n36056), .A1(n32630), .A2(n32629), .B0(conv_3[410]), 
        .B1(n32628), .Y(n32631) );
  NOR2X1 U20343 ( .A(n32627), .B(n32626), .Y(n32629) );
  AOI32XL U20344 ( .A0(n36056), .A1(n34142), .A2(n34141), .B0(conv_3[388]), 
        .B1(n34140), .Y(n34143) );
  NAND2XL U20345 ( .A(n34139), .B(n34138), .Y(n34141) );
  AOI2BB1XL U20346 ( .A0N(n34169), .A1N(n34168), .B0(n34167), .Y(n34170) );
  NOR2X1 U20347 ( .A(n34169), .B(n34166), .Y(n34165) );
  NOR2BXL U20348 ( .AN(n31642), .B(n31631), .Y(n31633) );
  NOR2X1 U20349 ( .A(n33833), .B(n33832), .Y(n33829) );
  NOR2X1 U20350 ( .A(n32128), .B(n32129), .Y(n31470) );
  NOR2X1 U20351 ( .A(n33752), .B(n33474), .Y(n33471) );
  NOR2X1 U20352 ( .A(n31480), .B(n31479), .Y(n31482) );
  AOI32XL U20353 ( .A0(n35748), .A1(n27592), .A2(n27591), .B0(n31957), .B1(
        n27592), .Y(n15519) );
  NOR2X1 U20354 ( .A(n35754), .B(n35753), .Y(n35755) );
  AOI32XL U20355 ( .A0(n36056), .A1(n34070), .A2(n34069), .B0(conv_3[328]), 
        .B1(n34068), .Y(n34071) );
  NAND2XL U20356 ( .A(n34067), .B(n34066), .Y(n34069) );
  NOR2X1 U20357 ( .A(n35740), .B(n35739), .Y(n35741) );
  AOI32XL U20358 ( .A0(n35743), .A1(n28761), .A2(n28760), .B0(n31908), .B1(
        n28761), .Y(n15532) );
  AOI32XL U20359 ( .A0(n36056), .A1(n34034), .A2(n34033), .B0(conv_3[313]), 
        .B1(n34032), .Y(n34035) );
  NAND2XL U20360 ( .A(n34031), .B(n34030), .Y(n34033) );
  AOI2BB1XL U20361 ( .A0N(n32540), .A1N(n35736), .B0(n32539), .Y(n32541) );
  NOR2X1 U20362 ( .A(n32540), .B(n32538), .Y(n32537) );
  AOI2BB1XL U20363 ( .A0N(n34483), .A1N(n35726), .B0(n34482), .Y(n34484) );
  NOR2X1 U20364 ( .A(n34483), .B(n34481), .Y(n34480) );
  AOI31XL U20365 ( .A0(n36056), .A1(n35728), .A2(n35727), .B0(n16653), .Y(
        n35729) );
  NOR2X1 U20366 ( .A(n32603), .B(n32601), .Y(n32600) );
  NOR2X1 U20367 ( .A(n31732), .B(n26331), .Y(n26330) );
  AOI32XL U20368 ( .A0(n36056), .A1(n34249), .A2(n34248), .B0(conv_3[245]), 
        .B1(n34247), .Y(n34250) );
  NOR2X1 U20369 ( .A(n34653), .B(n34651), .Y(n34650) );
  OAI2BB1XL U20370 ( .A0N(conv_3[221]), .A1N(n35670), .B0(n35669), .Y(n15597)
         );
  AOI31XL U20371 ( .A0(n36056), .A1(n35668), .A2(n35667), .B0(n16653), .Y(
        n35669) );
  NOR2X1 U20372 ( .A(n35660), .B(n32059), .Y(n32056) );
  AOI32XL U20373 ( .A0(n35665), .A1(n28835), .A2(n28834), .B0(n31530), .B1(
        n28835), .Y(n15601) );
  AOI31XL U20374 ( .A0(n36056), .A1(n31531), .A2(n28832), .B0(n16653), .Y(
        n28835) );
  AOI32XL U20375 ( .A0(n36056), .A1(n28830), .A2(n26528), .B0(conv_3[215]), 
        .B1(n26527), .Y(n26529) );
  NOR2X1 U20376 ( .A(n28829), .B(n28831), .Y(n26528) );
  AOI32XL U20377 ( .A0(n35646), .A1(n28840), .A2(n28839), .B0(n31847), .B1(
        n28840), .Y(n15609) );
  AOI31XL U20378 ( .A0(n36056), .A1(n31849), .A2(n28837), .B0(n16653), .Y(
        n28840) );
  NOR2X1 U20379 ( .A(n34660), .B(n34658), .Y(n34657) );
  OAI2BB1XL U20380 ( .A0N(conv_3[200]), .A1N(n35650), .B0(n35649), .Y(n15613)
         );
  AOI31XL U20381 ( .A0(n36056), .A1(n35648), .A2(n35647), .B0(n16653), .Y(
        n35649) );
  NOR2X1 U20382 ( .A(n31620), .B(n31621), .Y(n31604) );
  NOR2X1 U20383 ( .A(n34703), .B(n34702), .Y(n34705) );
  OAI32XL U20384 ( .A0(conv_3[193]), .A1(n32208), .A2(n32207), .B0(n32206), 
        .B1(n32205), .Y(n32210) );
  OAI2BB1XL U20385 ( .A0N(conv_3[172]), .A1N(n35634), .B0(n35633), .Y(n15631)
         );
  AOI31XL U20386 ( .A0(n36056), .A1(n35632), .A2(n35631), .B0(n16653), .Y(
        n35633) );
  NOR2X1 U20387 ( .A(n31585), .B(n31584), .Y(n31587) );
  NOR2X1 U20388 ( .A(n32285), .B(n32284), .Y(n32287) );
  AOI32XL U20389 ( .A0(n36056), .A1(n34754), .A2(n34753), .B0(conv_3[150]), 
        .B1(n34752), .Y(n34756) );
  NOR2X1 U20390 ( .A(n33971), .B(n33969), .Y(n33968) );
  NOR2X1 U20391 ( .A(n33466), .B(n33465), .Y(n33462) );
  NOR2X1 U20392 ( .A(n31714), .B(n31713), .Y(n31716) );
  AOI2BB1XL U20393 ( .A0N(n34400), .A1N(n34737), .B0(n34399), .Y(n34401) );
  NOR2X1 U20394 ( .A(n33709), .B(n33710), .Y(n31440) );
  NOR2X1 U20395 ( .A(n35622), .B(n33797), .Y(n33794) );
  NOR2X1 U20396 ( .A(n31399), .B(n31398), .Y(n31401) );
  AOI2BB1XL U20397 ( .A0N(n34201), .A1N(n34200), .B0(n34199), .Y(n34202) );
  NOR2X1 U20398 ( .A(n34201), .B(n34198), .Y(n34197) );
  NOR2X1 U20399 ( .A(n32640), .B(n32638), .Y(n32637) );
  AOI32XL U20400 ( .A0(n36056), .A1(n32669), .A2(n32668), .B0(conv_3[103]), 
        .B1(n32667), .Y(n32670) );
  OAI21XL U20401 ( .A0(n16654), .A1(n32668), .B0(n35618), .Y(n32667) );
  NAND2XL U20402 ( .A(n32666), .B(n32665), .Y(n32668) );
  AOI2BB1XL U20403 ( .A0N(n34192), .A1N(n35618), .B0(n34191), .Y(n34193) );
  NOR2X1 U20404 ( .A(n34192), .B(n34190), .Y(n34189) );
  AOI2BB1XL U20405 ( .A0N(n34184), .A1N(n35618), .B0(n34183), .Y(n34185) );
  NOR2X1 U20406 ( .A(n34184), .B(n34182), .Y(n34181) );
  AOI2BB1XL U20407 ( .A0N(n34186), .A1N(n32114), .B0(n32115), .Y(n31670) );
  NOR2X1 U20408 ( .A(n31680), .B(n31679), .Y(n31682) );
  AOI32XL U20409 ( .A0(n36056), .A1(n32573), .A2(n32572), .B0(conv_3[73]), 
        .B1(n32571), .Y(n32574) );
  OAI21XL U20410 ( .A0(n16654), .A1(n32572), .B0(n35598), .Y(n32571) );
  NAND2XL U20411 ( .A(n32570), .B(n32569), .Y(n32572) );
  AOI32XL U20412 ( .A0(n36056), .A1(n34160), .A2(n34159), .B0(conv_3[58]), 
        .B1(n34158), .Y(n34161) );
  AOI2BB1XL U20413 ( .A0N(n34393), .A1N(n34392), .B0(n34391), .Y(n34394) );
  NOR2X1 U20414 ( .A(n34393), .B(n34390), .Y(n34388) );
  AOI2BB1XL U20415 ( .A0N(n34375), .A1N(n34392), .B0(n34374), .Y(n34376) );
  NOR2X1 U20416 ( .A(n34375), .B(n34373), .Y(n34372) );
  AOI32XL U20417 ( .A0(n36056), .A1(n34414), .A2(n34413), .B0(conv_3[28]), 
        .B1(n34412), .Y(n34415) );
  AOI32XL U20418 ( .A0(n34383), .A1(n28642), .A2(n28641), .B0(n28640), .B1(
        n28642), .Y(n15736) );
  AOI2BB1XL U20419 ( .A0N(n34384), .A1N(n34383), .B0(n34382), .Y(n34385) );
  OAI211XL U20420 ( .A0(n34789), .A1(n33160), .B0(n33468), .C0(n33159), .Y(
        n15734) );
  AOI2BB2XL U20421 ( .B0(n36114), .B1(n36108), .A0N(filter_1_bias[0]), .A1N(
        n36114), .Y(n14733) );
  AOI2BB2XL U20422 ( .B0(n36107), .B1(n36106), .A0N(filter_3[1]), .A1N(n36107), 
        .Y(n14736) );
  AOI2BB2XL U20423 ( .B0(n36107), .B1(n36105), .A0N(filter_3[2]), .A1N(n36107), 
        .Y(n14737) );
  AOI2BB2XL U20424 ( .B0(n36107), .B1(n36104), .A0N(filter_3[3]), .A1N(n36107), 
        .Y(n14738) );
  AOI2BB2XL U20425 ( .B0(n36107), .B1(n36103), .A0N(filter_3[4]), .A1N(n36107), 
        .Y(n14739) );
  AOI2BB2XL U20426 ( .B0(n36107), .B1(n36102), .A0N(filter_3[5]), .A1N(n36107), 
        .Y(n14740) );
  AOI2BB2XL U20427 ( .B0(n36107), .B1(n36101), .A0N(filter_3[0]), .A1N(n36107), 
        .Y(n14741) );
  AOI2BB2XL U20428 ( .B0(n36100), .B1(n36099), .A0N(filter_2[1]), .A1N(n20603), 
        .Y(n14790) );
  AOI2BB2XL U20429 ( .B0(n36100), .B1(n36098), .A0N(filter_2[2]), .A1N(n20603), 
        .Y(n14791) );
  AOI2BB2XL U20430 ( .B0(n36100), .B1(n36097), .A0N(filter_2[3]), .A1N(n20603), 
        .Y(n14792) );
  AOI2BB2XL U20431 ( .B0(n36100), .B1(n36096), .A0N(filter_2[4]), .A1N(n20603), 
        .Y(n14793) );
  AOI2BB2XL U20432 ( .B0(n36100), .B1(n36095), .A0N(filter_2[5]), .A1N(n20603), 
        .Y(n14794) );
  AOI2BB2XL U20433 ( .B0(n36100), .B1(n36094), .A0N(filter_2[0]), .A1N(n20603), 
        .Y(n14795) );
  OAI31XL U20434 ( .A0(n35255), .A1(n19187), .A2(n19224), .B0(n19186), .Y(
        n16642) );
  AOI22XL U20435 ( .A0(N18014), .A1(n19222), .B0(n35256), .B1(N29499), .Y(
        n19186) );
  AOI2BB2XL U20436 ( .B0(n22896), .B1(n35254), .A0N(pixel[0]), .A1N(n22896), 
        .Y(N17494) );
  AOI211XL U20437 ( .A0(n18773), .A1(counter[5]), .B0(n19242), .C0(n26848), 
        .Y(N30144) );
  OAI31X1 U20438 ( .A0(n18182), .A1(n18165), .A2(n18164), .B0(n36247), .Y(
        n18166) );
  AOI211XL U20439 ( .A0(n18191), .A1(n19004), .B0(cs[1]), .C0(n18175), .Y(
        n18165) );
  OAI32XL U20440 ( .A0(n18176), .A1(n18190), .A2(n18163), .B0(cs[0]), .B1(
        n18162), .Y(n18164) );
  NOR2X4 U20441 ( .A(N17708), .B(n18516), .Y(n22347) );
  AOI221X2 U20442 ( .A0(n19695), .A1(n18106), .B0(n18107), .B1(n19697), .C0(
        n19696), .Y(n18154) );
  AND2X4 U20443 ( .A(ns[0]), .B(n19183), .Y(n36056) );
  OAI21X2 U20444 ( .A0(n18184), .A1(n18187), .B0(n18166), .Y(ns[0]) );
  OAI211XL U20445 ( .A0(n33443), .A1(n33442), .B0(n34544), .C0(n33441), .Y(
        n16434) );
  NAND2XL U20446 ( .A(conv_1[29]), .B(n33440), .Y(n33439) );
  AOI22XL U20447 ( .A0(conv_1[28]), .A1(n33438), .B0(n33437), .B1(n33436), .Y(
        n33440) );
  AOI221X1 U20448 ( .A0(n19636), .A1(n17962), .B0(n17963), .B1(n19638), .C0(
        n19637), .Y(n18003) );
  NAND2XL U20449 ( .A(n30414), .B(conv_2[167]), .Y(n30413) );
  NOR2X4 U20450 ( .A(n21358), .B(n18516), .Y(n16723) );
  INVX4 U20451 ( .A(n16723), .Y(n22716) );
  INVX4 U20452 ( .A(n18286), .Y(n22770) );
  ADDFHX1 U20453 ( .A(DP_OP_5167J1_123_9881_n22), .B(DP_OP_5167J1_123_9881_n27), .CI(n22196), .CO(n25242), .S(n20724) );
  OAI31XL U20454 ( .A0(n17439), .A1(n17438), .A2(n17437), .B0(n19182), .Y(
        n17440) );
  OAI2BB1X2 U20455 ( .A0N(conv_3[9]), .A1N(n31159), .B0(n24373), .Y(n28637) );
  OAI2BB1XL U20456 ( .A0N(conv_3[2]), .A1N(n30786), .B0(n23756), .Y(n24330) );
  NAND2X2 U20457 ( .A(n22896), .B(filter_3_bias[5]), .Y(n35588) );
  NOR2X4 U20458 ( .A(n36244), .B(n28292), .Y(n22369) );
  XOR2X1 U20459 ( .A(n33558), .B(n33557), .Y(n33559) );
  NAND2X2 U20460 ( .A(N18014), .B(n28467), .Y(n16701) );
  OAI2BB2XL U20461 ( .B0(n33410), .B1(n33409), .A0N(n33410), .A1N(n33409), .Y(
        n33411) );
  XOR2X1 U20462 ( .A(n33408), .B(n33407), .Y(n33409) );
  NAND2XL U20463 ( .A(n33980), .B(n35970), .Y(n34022) );
  AOI2BB1XL U20464 ( .A0N(conv_1[96]), .A1N(n26789), .B0(n31334), .Y(n26807)
         );
  INVX12 U20465 ( .A(n18208), .Y(n35236) );
  NOR2X2 U20466 ( .A(n19221), .B(n28467), .Y(n16700) );
  AOI2BB1X2 U20467 ( .A0N(conv_1[377]), .A1N(n23723), .B0(n23724), .Y(n23193)
         );
  AND2X2 U20468 ( .A(n19148), .B(n19149), .Y(n23723) );
  OAI211XL U20469 ( .A0(n33853), .A1(n33152), .B0(n34281), .C0(n33151), .Y(
        n16074) );
  NAND2XL U20470 ( .A(conv_1[389]), .B(n33150), .Y(n33149) );
  AOI22XL U20471 ( .A0(conv_1[388]), .A1(n33148), .B0(n33147), .B1(n33146), 
        .Y(n33150) );
  ADDFHX1 U20472 ( .A(conv_2[171]), .B(n29831), .CI(n30968), .CO(n29846), .S(
        n30970) );
  AOI2BB1XL U20473 ( .A0N(conv_2[170]), .A1N(n29840), .B0(n29839), .Y(n30968)
         );
  AOI22XL U20474 ( .A0(conv_2[178]), .A1(n34594), .B0(n34593), .B1(n34592), 
        .Y(n34596) );
  NOR3X2 U20475 ( .A(n33989), .B(n22257), .C(n34434), .Y(n34431) );
  NAND2XL U20476 ( .A(conv_3[479]), .B(n32187), .Y(n32186) );
  AOI22XL U20477 ( .A0(conv_3[478]), .A1(n32322), .B0(n32321), .B1(n32326), 
        .Y(n32187) );
  INVX3 U20478 ( .A(n22362), .Y(n25123) );
  NAND2X4 U20479 ( .A(n19242), .B(n19183), .Y(n23672) );
  AND2X2 U20480 ( .A(n36244), .B(n36245), .Y(n22362) );
  AOI211X2 U20481 ( .A0(counter[3]), .A1(filter_3[50]), .B0(n18996), .C0(
        n18995), .Y(n18997) );
  INVXL U20482 ( .A(n18856), .Y(n33442) );
  NOR2X2 U20483 ( .A(n19183), .B(n29676), .Y(n18856) );
  INVXL U20484 ( .A(n18856), .Y(n34789) );
  INVXL U20485 ( .A(n18856), .Y(n34520) );
  INVXL U20486 ( .A(n18856), .Y(n34676) );
  NOR2X1 U20487 ( .A(n16721), .B(n18196), .Y(n18197) );
  INVX2 U20488 ( .A(n36244), .Y(n16721) );
  NOR2X2 U20489 ( .A(n36245), .B(n18239), .Y(n21954) );
  BUFX8 U20490 ( .A(N17785), .Y(n36245) );
  BUFX4 U20491 ( .A(n16702), .Y(n28292) );
  INVX2 U20492 ( .A(n22770), .Y(n19401) );
  INVX2 U20493 ( .A(n16700), .Y(n35135) );
  INVXL U20494 ( .A(n16700), .Y(n35241) );
  NOR2X2 U20495 ( .A(n18815), .B(n16701), .Y(n26263) );
  INVXL U20496 ( .A(n26470), .Y(n26479) );
  INVXL U20497 ( .A(n35588), .Y(n31384) );
  INVX2 U20498 ( .A(n16653), .Y(n33468) );
  INVX2 U20499 ( .A(n35159), .Y(n16755) );
  INVX2 U20500 ( .A(n34981), .Y(n28414) );
  INVXL U20501 ( .A(n16746), .Y(n34981) );
  INVX2 U20502 ( .A(n26621), .Y(n28324) );
  INVX2 U20503 ( .A(n28556), .Y(n28577) );
  INVXL U20504 ( .A(n16673), .Y(n24039) );
  INVX2 U20505 ( .A(n16715), .Y(n18810) );
  INVX2 U20506 ( .A(n16715), .Y(n25289) );
  INVX2 U20507 ( .A(n25289), .Y(n22612) );
  INVXL U20508 ( .A(n16668), .Y(n18658) );
  INVX2 U20509 ( .A(n18239), .Y(n22616) );
  INVX2 U20510 ( .A(n22759), .Y(n22717) );
  INVXL U20511 ( .A(n25299), .Y(n22550) );
  NOR2X2 U20512 ( .A(N17708), .B(n35269), .Y(n22368) );
  INVX2 U20513 ( .A(n19401), .Y(n20978) );
  INVX2 U20514 ( .A(n19902), .Y(n25306) );
  INVX2 U20515 ( .A(n19902), .Y(n22762) );
  INVX2 U20516 ( .A(n16706), .Y(n19416) );
  INVX2 U20517 ( .A(n28414), .Y(n28575) );
  NAND2X1 U20518 ( .A(n36245), .B(n16755), .Y(n28349) );
  INVXL U20519 ( .A(n21762), .Y(n21556) );
  INVXL U20520 ( .A(n21887), .Y(n21810) );
  INVX2 U20521 ( .A(n26479), .Y(n35130) );
  INVX2 U20522 ( .A(n34827), .Y(n26575) );
  INVX2 U20523 ( .A(n35241), .Y(n28465) );
  INVX2 U20524 ( .A(n18197), .Y(n35198) );
  INVXL U20525 ( .A(n28479), .Y(n34992) );
  NOR2X1 U20526 ( .A(n18815), .B(n35159), .Y(n16745) );
  INVX2 U20527 ( .A(n26853), .Y(n32491) );
  INVXL U20528 ( .A(n26853), .Y(n31071) );
  INVXL U20529 ( .A(n26853), .Y(n26906) );
  INVXL U20530 ( .A(n26853), .Y(n31077) );
  INVX2 U20531 ( .A(n31077), .Y(n26910) );
  INVX2 U20532 ( .A(n16651), .Y(n34735) );
  INVX2 U20533 ( .A(n16651), .Y(n33815) );
  INVX2 U20534 ( .A(n16651), .Y(n34669) );
  NOR2X2 U20535 ( .A(n36249), .B(n19610), .Y(n16674) );
  INVX2 U20536 ( .A(n20603), .Y(n22105) );
  INVXL U20537 ( .A(n33912), .Y(n34389) );
  INVX2 U20538 ( .A(n16658), .Y(n35336) );
  INVXL U20539 ( .A(n36042), .Y(n33157) );
  INVXL U20540 ( .A(n36042), .Y(n24378) );
  INVXL U20541 ( .A(n33912), .Y(n36009) );
  INVX2 U20542 ( .A(n36001), .Y(n33778) );
  INVXL U20543 ( .A(n36001), .Y(n34666) );
  INVXL U20544 ( .A(n36001), .Y(n27932) );
  INVXL U20545 ( .A(n36001), .Y(n33712) );
  INVXL U20546 ( .A(n36042), .Y(n24499) );
  INVXL U20547 ( .A(n36001), .Y(n32660) );
  INVX2 U20548 ( .A(n16658), .Y(n36020) );
  INVXL U20549 ( .A(n36042), .Y(n28751) );
  INVXL U20550 ( .A(n16656), .Y(n35419) );
  INVXL U20551 ( .A(n36001), .Y(n32052) );
  INVXL U20552 ( .A(n36001), .Y(n30090) );
  INVXL U20553 ( .A(n36001), .Y(n31735) );
  INVX2 U20554 ( .A(n36056), .Y(n36042) );
  INVXL U20555 ( .A(n17969), .Y(n19698) );
  AOI222XL U20556 ( .A0(counter[1]), .A1(affine_1[20]), .B0(n17988), .B1(
        affine_1[10]), .C0(n19228), .C1(affine_1[0]), .Y(n17969) );
  INVXL U20557 ( .A(n19698), .Y(n19652) );
  INVX2 U20558 ( .A(n20608), .Y(n28249) );
  INVX2 U20559 ( .A(n28249), .Y(n36120) );
  INVXL U20560 ( .A(n33403), .Y(n24909) );
  AOI211X2 U20561 ( .A0(counter[3]), .A1(filter_1[50]), .B0(n18834), .C0(
        n18833), .Y(n33403) );
  INVXL U20562 ( .A(n17936), .Y(n24570) );
  NOR2X1 U20563 ( .A(n16715), .B(n26274), .Y(n17866) );
  NOR2X1 U20564 ( .A(n19902), .B(n23186), .Y(n19904) );
  INVXL U20565 ( .A(n26027), .Y(n21925) );
  INVXL U20566 ( .A(n35089), .Y(n26216) );
  INVXL U20567 ( .A(n18109), .Y(n18115) );
  INVXL U20568 ( .A(n25515), .Y(n24730) );
  INVXL U20569 ( .A(n19427), .Y(n21371) );
  INVXL U20570 ( .A(n28321), .Y(n35066) );
  OAI2BB1X1 U20571 ( .A0N(weight_2[51]), .A1N(n18049), .B0(n18036), .Y(n19614)
         );
  INVXL U20572 ( .A(n17949), .Y(n18141) );
  INVXL U20573 ( .A(n28421), .Y(n26633) );
  INVXL U20574 ( .A(n26083), .Y(n22027) );
  INVXL U20575 ( .A(n25726), .Y(n35061) );
  INVXL U20576 ( .A(n35184), .Y(n35207) );
  INVXL U20577 ( .A(n18106), .Y(n19697) );
  INVXL U20578 ( .A(n30525), .Y(n23060) );
  INVXL U20579 ( .A(n21464), .Y(n21311) );
  INVXL U20580 ( .A(n35104), .Y(n24828) );
  INVXL U20581 ( .A(n20580), .Y(n20586) );
  INVX2 U20582 ( .A(n17026), .Y(n19007) );
  XOR2XL U20583 ( .A(affine_1[14]), .B(n17505), .Y(DP_OP_5167J1_123_9881_n40)
         );
  XOR2XL U20584 ( .A(affine_2[10]), .B(n18155), .Y(DP_OP_5171J1_127_4278_n36)
         );
  INVXL U20585 ( .A(n18010), .Y(n19630) );
  NOR2X1 U20586 ( .A(n27214), .B(n27213), .Y(n27215) );
  INVXL U20587 ( .A(n20207), .Y(n21479) );
  INVXL U20588 ( .A(n20755), .Y(n18204) );
  INVXL U20589 ( .A(n21004), .Y(n21678) );
  AOI222XL U20590 ( .A0(n27386), .A1(n27387), .B0(n27386), .B1(conv_1[514]), 
        .C0(n27387), .C1(conv_1[514]), .Y(n24912) );
  NOR2X2 U20591 ( .A(n16721), .B(n17170), .Y(n22015) );
  ADDFXL U20592 ( .A(n20622), .B(n20621), .CI(n20620), .CO(n20695), .S(n20680)
         );
  NOR2X1 U20593 ( .A(n23822), .B(n23824), .Y(n23820) );
  NOR2X1 U20594 ( .A(n23888), .B(n23886), .Y(n23884) );
  INVXL U20595 ( .A(n25119), .Y(n25496) );
  INVX4 U20596 ( .A(n35239), .Y(n35195) );
  INVXL U20597 ( .A(n18997), .Y(n27619) );
  INVXL U20598 ( .A(n24956), .Y(n24962) );
  NOR2X1 U20599 ( .A(n22220), .B(n26148), .Y(n23696) );
  INVXL U20600 ( .A(n21458), .Y(n21463) );
  AOI221XL U20601 ( .A0(n22705), .A1(n22799), .B0(n22704), .B1(n22799), .C0(
        n22703), .Y(n22794) );
  INVXL U20602 ( .A(n34768), .Y(n35499) );
  INVXL U20603 ( .A(n28821), .Y(n35434) );
  INVXL U20604 ( .A(n34259), .Y(n29382) );
  INVXL U20605 ( .A(n34019), .Y(n27764) );
  INVXL U20606 ( .A(n33780), .Y(n31517) );
  INVXL U20607 ( .A(n34525), .Y(n34522) );
  INVXL U20608 ( .A(n32618), .Y(n32599) );
  INVXL U20609 ( .A(n23016), .Y(n23789) );
  INVXL U20610 ( .A(n34379), .Y(n32996) );
  ADDFXL U20611 ( .A(conv_2[107]), .B(n25676), .CI(n25675), .CO(n27140), .S(
        n23576) );
  XOR2XL U20612 ( .A(n30806), .B(n30805), .Y(n30808) );
  ADDFXL U20613 ( .A(conv_3[62]), .B(n24237), .CI(n24236), .CO(n23897), .S(
        n24238) );
  ADDFXL U20614 ( .A(conv_1[153]), .B(n24283), .CI(n24282), .CO(n24009), .S(
        n24284) );
  XOR2XL U20615 ( .A(n23234), .B(n23233), .Y(n23236) );
  AOI222XL U20616 ( .A0(n20098), .A1(n20097), .B0(n20098), .B1(n20096), .C0(
        n20097), .C1(n20095), .Y(n20099) );
  INVXL U20617 ( .A(n34852), .Y(n26381) );
  INVXL U20618 ( .A(n33424), .Y(n33422) );
  NAND4X1 U20619 ( .A(n22854), .B(n22853), .C(n22852), .D(n22851), .Y(n34717)
         );
  ADDFXL U20620 ( .A(conv_1[8]), .B(n27278), .CI(n22383), .CO(n24537), .S(
        n22384) );
  AOI222XL U20621 ( .A0(n22046), .A1(n22045), .B0(n22046), .B1(n22044), .C0(
        n22045), .C1(n22043), .Y(n22047) );
  ADDFXL U20622 ( .A(conv_2[367]), .B(n34570), .CI(n24454), .CO(n29507), .S(
        n24456) );
  ADDFXL U20623 ( .A(conv_2[321]), .B(n35982), .CI(n26352), .CO(n35983), .S(
        n23107) );
  NOR2X1 U20624 ( .A(conv_2[72]), .B(n33732), .Y(n33733) );
  INVXL U20625 ( .A(n33620), .Y(n28673) );
  AOI222XL U20626 ( .A0(n35226), .A1(n35225), .B0(n35226), .B1(n35224), .C0(
        n35225), .C1(n35223), .Y(n35228) );
  ADDFXL U20627 ( .A(conv_3[515]), .B(n31180), .CI(n24478), .CO(n31173), .S(
        n24460) );
  ADDFXL U20628 ( .A(conv_3[383]), .B(n34164), .CI(n32525), .CO(n31502), .S(
        n32526) );
  INVXL U20629 ( .A(n33842), .Y(n33281) );
  INVXL U20630 ( .A(n19108), .Y(n33867) );
  NOR2X1 U20631 ( .A(conv_3[129]), .B(n28953), .Y(n31438) );
  INVXL U20632 ( .A(in_data[9]), .Y(n20167) );
  NAND2X1 U20633 ( .A(n36123), .B(n30349), .Y(n20416) );
  INVXL U20634 ( .A(n23663), .Y(n33427) );
  INVXL U20635 ( .A(n35510), .Y(n35504) );
  INVXL U20636 ( .A(n33649), .Y(n35477) );
  INVXL U20637 ( .A(n22318), .Y(n22317) );
  AOI32XL U20638 ( .A0(n36056), .A1(n29251), .A2(n27968), .B0(conv_1[283]), 
        .B1(n27967), .Y(n27969) );
  AOI32XL U20639 ( .A0(n36056), .A1(n26496), .A2(n26495), .B0(conv_1[251]), 
        .B1(n26494), .Y(n26497) );
  AOI32XL U20640 ( .A0(n36056), .A1(n33846), .A2(n33486), .B0(conv_1[238]), 
        .B1(n33485), .Y(n33487) );
  INVXL U20641 ( .A(n23915), .Y(n35346) );
  INVXL U20642 ( .A(n35341), .Y(n34271) );
  AOI31XL U20643 ( .A0(n36056), .A1(n36055), .A2(n36054), .B0(n16651), .Y(
        n36057) );
  INVXL U20644 ( .A(n18856), .Y(n33853) );
  INVXL U20645 ( .A(n24303), .Y(n36003) );
  INVXL U20646 ( .A(n35952), .Y(n30994) );
  AOI31XL U20647 ( .A0(n36056), .A1(n35937), .A2(n35936), .B0(n16651), .Y(
        n35938) );
  INVXL U20648 ( .A(n33765), .Y(n35934) );
  INVXL U20649 ( .A(n24358), .Y(n34631) );
  INVXL U20650 ( .A(n33774), .Y(n35805) );
  INVXL U20651 ( .A(n32546), .Y(n34227) );
  AOI31XL U20652 ( .A0(n36056), .A1(n35709), .A2(n35708), .B0(n16653), .Y(
        n35710) );
  AOI32XL U20653 ( .A0(n36056), .A1(n33898), .A2(n33882), .B0(conv_3[238]), 
        .B1(n33881), .Y(n33883) );
  INVXL U20654 ( .A(n33444), .Y(n35594) );
  NAND2BX1 U20655 ( .AN(n30350), .B(n30349), .Y(n30392) );
  OAI21XL U20656 ( .A0(in_data[8]), .A1(in_data[7]), .B0(n20168), .Y(n36124)
         );
  AOI22XL U20657 ( .A0(counter[1]), .A1(pool[130]), .B0(counter[0]), .B1(
        pool[125]), .Y(n16699) );
  INVXL U20658 ( .A(n19005), .Y(n17028) );
  NOR2X2 U20659 ( .A(counter[1]), .B(counter[0]), .Y(n19228) );
  INVXL U20660 ( .A(n17027), .Y(n16987) );
  NAND2XL U20661 ( .A(counter[3]), .B(n16987), .Y(n17017) );
  AOI22XL U20662 ( .A0(pool[50]), .A1(n17011), .B0(pool[40]), .B1(n17010), .Y(
        n16698) );
  INVXL U20663 ( .A(n18156), .Y(n17006) );
  NAND2X1 U20664 ( .A(counter[2]), .B(n19228), .Y(n17026) );
  AOI22XL U20665 ( .A0(n19004), .A1(pool[25]), .B0(n19007), .B1(pool[20]), .Y(
        n16680) );
  AOI22XL U20666 ( .A0(n19009), .A1(pool[15]), .B0(n19006), .B1(pool[5]), .Y(
        n16679) );
  AOI22XL U20667 ( .A0(n19005), .A1(pool[10]), .B0(n16987), .B1(pool[0]), .Y(
        n16678) );
  AOI22XL U20668 ( .A0(n19008), .A1(pool[35]), .B0(n16676), .B1(pool[30]), .Y(
        n16677) );
  NAND4XL U20669 ( .A(n16680), .B(n16679), .C(n16678), .D(n16677), .Y(n16696)
         );
  INVXL U20670 ( .A(pool[80]), .Y(n34922) );
  AOI22XL U20671 ( .A0(n19007), .A1(pool[100]), .B0(n19005), .B1(pool[90]), 
        .Y(n16682) );
  NAND2XL U20672 ( .A(n19006), .B(pool[85]), .Y(n16681) );
  OAI211XL U20673 ( .A0(n34922), .A1(n17027), .B0(n16682), .C0(n16681), .Y(
        n16689) );
  INVXL U20674 ( .A(n17017), .Y(n16683) );
  AOI22XL U20675 ( .A0(n19008), .A1(pool[115]), .B0(pool[120]), .B1(n16683), 
        .Y(n16684) );
  OAI2BB1XL U20676 ( .A0N(n19004), .A1N(pool[105]), .B0(n16684), .Y(n16688) );
  AOI22XL U20677 ( .A0(n19009), .A1(pool[95]), .B0(n16676), .B1(pool[110]), 
        .Y(n16686) );
  OAI31XL U20678 ( .A0(pool[60]), .A1(pool[120]), .A2(pool[100]), .B0(n19228), 
        .Y(n16685) );
  INVXL U20679 ( .A(n20363), .Y(n18170) );
  AOI32XL U20680 ( .A0(n16699), .A1(n16686), .A2(n16685), .B0(n18170), .B1(
        n16686), .Y(n16687) );
  AOI211XL U20681 ( .A0(n19247), .A1(n16689), .B0(n16688), .C0(n16687), .Y(
        n16694) );
  AOI22XL U20682 ( .A0(n18159), .A1(pool[45]), .B0(pool[60]), .B1(n17038), .Y(
        n16693) );
  AOI22XL U20683 ( .A0(n19009), .A1(pool[55]), .B0(n16676), .B1(pool[70]), .Y(
        n16691) );
  AOI22XL U20684 ( .A0(n19008), .A1(pool[75]), .B0(n19004), .B1(pool[65]), .Y(
        n16690) );
  OAI2BB1XL U20685 ( .A0N(n16691), .A1N(n16690), .B0(counter[3]), .Y(n16692)
         );
  OAI211XL U20686 ( .A0(n16694), .A1(n20600), .B0(n16693), .C0(n16692), .Y(
        n16695) );
  AOI21XL U20687 ( .A0(n17006), .A1(n16696), .B0(n16695), .Y(n16697) );
  NOR2X4 U20688 ( .A(n19855), .B(n21830), .Y(n19098) );
  INVX8 U20689 ( .A(N18471), .Y(n28467) );
  INVXL U20690 ( .A(n17800), .Y(n16951) );
  INVXL U20691 ( .A(weight_1[454]), .Y(n32386) );
  INVX4 U20692 ( .A(n22347), .Y(n18286) );
  NOR2X1 U20693 ( .A(n26575), .B(n19182), .Y(n17169) );
  INVXL U20694 ( .A(weight_1[448]), .Y(n32385) );
  INVXL U20695 ( .A(n17169), .Y(n16707) );
  OAI22XL U20696 ( .A0(n32386), .A1(n17746), .B0(n32385), .B1(n17690), .Y(
        n16705) );
  INVXL U20697 ( .A(weight_1[478]), .Y(n32759) );
  INVX2 U20698 ( .A(n36245), .Y(n16702) );
  NOR2X4 U20699 ( .A(n26374), .B(n18286), .Y(n19099) );
  INVXL U20700 ( .A(n17842), .Y(n17694) );
  INVXL U20701 ( .A(weight_1[472]), .Y(n32760) );
  NOR2X1 U20702 ( .A(n28292), .B(n18239), .Y(n16703) );
  NAND2X1 U20703 ( .A(n34827), .B(n19475), .Y(n21731) );
  NAND2XL U20704 ( .A(n21749), .B(cursor[6]), .Y(n17846) );
  OAI22XL U20705 ( .A0(n32759), .A1(n17694), .B0(n32760), .B1(n17846), .Y(
        n16704) );
  AOI211XL U20706 ( .A0(weight_1[10]), .A1(n17444), .B0(n16705), .C0(n16704), 
        .Y(n16777) );
  NAND2XL U20707 ( .A(n21887), .B(n17169), .Y(n17747) );
  INVX4 U20708 ( .A(N17708), .Y(n21358) );
  AOI22XL U20709 ( .A0(weight_1[466]), .A1(n17852), .B0(weight_1[460]), .B1(
        n17753), .Y(n16776) );
  NAND2XL U20710 ( .A(n34827), .B(n21831), .Y(n20491) );
  AOI2BB1XL U20711 ( .A0N(n17923), .A1N(n28467), .B0(n22011), .Y(n17144) );
  AOI22XL U20712 ( .A0(n22021), .A1(weight_1[412]), .B0(n16734), .B1(
        weight_1[406]), .Y(n16713) );
  AOI22XL U20713 ( .A0(n19098), .A1(weight_1[442]), .B0(n19099), .B1(
        weight_1[430]), .Y(n16712) );
  AOI22XL U20714 ( .A0(n19097), .A1(weight_1[436]), .B0(n21887), .B1(
        weight_1[418]), .Y(n16711) );
  AOI22XL U20715 ( .A0(n19475), .A1(weight_1[424]), .B0(n21954), .B1(
        weight_1[400]), .Y(n16710) );
  NAND4XL U20716 ( .A(n16713), .B(n16712), .C(n16711), .D(n16710), .Y(n16714)
         );
  AOI22XL U20717 ( .A0(weight_1[484]), .A1(n17068), .B0(n17166), .B1(n16714), 
        .Y(n16775) );
  INVXL U20718 ( .A(weight_1[196]), .Y(n32959) );
  INVX2 U20719 ( .A(n16715), .Y(n16716) );
  INVXL U20720 ( .A(weight_1[394]), .Y(n32452) );
  INVXL U20721 ( .A(n17813), .Y(n17391) );
  INVXL U20722 ( .A(weight_1[4]), .Y(n32910) );
  OAI22XL U20723 ( .A0(n32452), .A1(n17391), .B0(n32910), .B1(n17188), .Y(
        n16772) );
  NOR2X4 U20724 ( .A(N18014), .B(n28467), .Y(n26470) );
  NOR2X1 U20725 ( .A(n26479), .B(n16721), .Y(n23055) );
  INVXL U20726 ( .A(n23055), .Y(n16760) );
  AOI22XL U20727 ( .A0(n21766), .A1(weight_1[322]), .B0(weight_1[394]), .B1(
        n17800), .Y(n16720) );
  AOI22XL U20728 ( .A0(weight_1[304]), .A1(n17798), .B0(weight_1[106]), .B1(
        n17885), .Y(n16719) );
  NOR2X4 U20729 ( .A(n36244), .B(n36245), .Y(n22370) );
  NOR2X2 U20730 ( .A(n22717), .B(n34981), .Y(n21762) );
  NOR2X2 U20731 ( .A(n26479), .B(n18815), .Y(n26276) );
  INVX2 U20732 ( .A(n26276), .Y(n26162) );
  NOR2X1 U20733 ( .A(n18286), .B(n26162), .Y(n17894) );
  AOI22XL U20734 ( .A0(n21762), .A1(weight_1[16]), .B0(weight_1[142]), .B1(
        n17894), .Y(n16718) );
  AOI22XL U20735 ( .A0(weight_1[292]), .A1(n17900), .B0(weight_1[166]), .B1(
        n17863), .Y(n16717) );
  NAND4XL U20736 ( .A(n16720), .B(n16719), .C(n16718), .D(n16717), .Y(n16743)
         );
  NOR2X1 U20737 ( .A(N18014), .B(n36245), .Y(n16722) );
  NAND2X1 U20738 ( .A(n16723), .B(n28290), .Y(n18109) );
  AOI22XL U20739 ( .A0(weight_1[226]), .A1(n17878), .B0(weight_1[76]), .B1(
        n17865), .Y(n16729) );
  INVX2 U20740 ( .A(n26085), .Y(n26059) );
  NAND2X1 U20741 ( .A(n22770), .B(n28290), .Y(n18117) );
  AOI22XL U20742 ( .A0(n26059), .A1(weight_1[334]), .B0(weight_1[214]), .B1(
        n17898), .Y(n16728) );
  AOI22XL U20743 ( .A0(weight_1[184]), .A1(n16724), .B0(weight_1[52]), .B1(
        n17803), .Y(n16727) );
  NOR2X1 U20744 ( .A(n16715), .B(n16661), .Y(n17897) );
  AOI22XL U20745 ( .A0(weight_1[124]), .A1(n17792), .B0(weight_1[100]), .B1(
        n17897), .Y(n16726) );
  NAND4XL U20746 ( .A(n16729), .B(n16728), .C(n16727), .D(n16726), .Y(n16742)
         );
  AOI22XL U20747 ( .A0(weight_1[382]), .A1(n17810), .B0(weight_1[376]), .B1(
        n17809), .Y(n16733) );
  AOI22XL U20748 ( .A0(weight_1[370]), .A1(n17825), .B0(weight_1[154]), .B1(
        n17822), .Y(n16732) );
  INVX4 U20749 ( .A(n35130), .Y(n34989) );
  NOR2X1 U20750 ( .A(n34989), .B(n22018), .Y(n17814) );
  AOI22XL U20751 ( .A0(weight_1[340]), .A1(n17814), .B0(weight_1[244]), .B1(
        n17815), .Y(n16731) );
  AOI22XL U20752 ( .A0(weight_1[352]), .A1(n17812), .B0(weight_1[202]), .B1(
        n17813), .Y(n16730) );
  NAND4XL U20753 ( .A(n16733), .B(n16732), .C(n16731), .D(n16730), .Y(n16741)
         );
  NAND2X2 U20754 ( .A(n19099), .B(n19221), .Y(n18120) );
  AOI22XL U20755 ( .A0(weight_1[238]), .A1(n17824), .B0(weight_1[70]), .B1(
        n17883), .Y(n16739) );
  AOI22XL U20756 ( .A0(weight_1[364]), .A1(n17827), .B0(weight_1[358]), .B1(
        n17816), .Y(n16738) );
  AOI22XL U20757 ( .A0(weight_1[388]), .A1(n17821), .B0(weight_1[346]), .B1(
        n17823), .Y(n16737) );
  NAND2XL U20758 ( .A(n19475), .B(n19221), .Y(n16735) );
  AOI22XL U20759 ( .A0(weight_1[298]), .A1(n17826), .B0(weight_1[232]), .B1(
        n17811), .Y(n16736) );
  NAND4XL U20760 ( .A(n16739), .B(n16738), .C(n16737), .D(n16736), .Y(n16740)
         );
  NOR4XL U20761 ( .A(n16743), .B(n16742), .C(n16741), .D(n16740), .Y(n16770)
         );
  AOI22XL U20762 ( .A0(weight_1[256]), .A1(n17896), .B0(weight_1[208]), .B1(
        n17884), .Y(n16750) );
  AOI22XL U20763 ( .A0(weight_1[268]), .A1(n17788), .B0(weight_1[64]), .B1(
        n17791), .Y(n16749) );
  INVX2 U20764 ( .A(n22030), .Y(n16744) );
  AOI22XL U20765 ( .A0(n16744), .A1(weight_1[88]), .B0(weight_1[40]), .B1(
        n17867), .Y(n16748) );
  NAND2XL U20766 ( .A(n23055), .B(n19475), .Y(n26029) );
  AOI22XL U20767 ( .A0(n26082), .A1(weight_1[328]), .B0(n21764), .B1(
        weight_1[22]), .Y(n16747) );
  NAND4XL U20768 ( .A(n16750), .B(n16749), .C(n16748), .D(n16747), .Y(n16768)
         );
  INVXL U20769 ( .A(n19099), .Y(n17173) );
  AOI22XL U20770 ( .A0(weight_1[286]), .A1(n17802), .B0(weight_1[58]), .B1(
        n17789), .Y(n16754) );
  AOI22XL U20771 ( .A0(n21748), .A1(weight_1[316]), .B0(weight_1[196]), .B1(
        n17866), .Y(n16753) );
  INVXL U20772 ( .A(n19475), .Y(n17165) );
  AOI22XL U20773 ( .A0(weight_1[280]), .A1(n17877), .B0(weight_1[46]), .B1(
        n17874), .Y(n16752) );
  AOI22XL U20774 ( .A0(weight_1[262]), .A1(n17886), .B0(weight_1[28]), .B1(
        n17893), .Y(n16751) );
  NAND4XL U20775 ( .A(n16754), .B(n16753), .C(n16752), .D(n16751), .Y(n16767)
         );
  NOR2X1 U20776 ( .A(n22717), .B(n26162), .Y(n17895) );
  AOI22XL U20777 ( .A0(weight_1[160]), .A1(n17868), .B0(weight_1[136]), .B1(
        n17895), .Y(n16759) );
  AOI22XL U20778 ( .A0(weight_1[250]), .A1(n17797), .B0(weight_1[178]), .B1(
        n17899), .Y(n16758) );
  AOI22XL U20779 ( .A0(weight_1[130]), .A1(n17801), .B0(weight_1[34]), .B1(
        n17873), .Y(n16757) );
  AOI22XL U20780 ( .A0(weight_1[172]), .A1(n17888), .B0(weight_1[112]), .B1(
        n17887), .Y(n16756) );
  NAND4XL U20781 ( .A(n16759), .B(n16758), .C(n16757), .D(n16756), .Y(n16766)
         );
  AOI22XL U20782 ( .A0(weight_1[274]), .A1(n17864), .B0(weight_1[118]), .B1(
        n17876), .Y(n16764) );
  AOI22XL U20783 ( .A0(weight_1[220]), .A1(n17804), .B0(weight_1[82]), .B1(
        n17799), .Y(n16763) );
  AOI22XL U20784 ( .A0(n21999), .A1(weight_1[94]), .B0(weight_1[148]), .B1(
        n17875), .Y(n16762) );
  AOI22XL U20785 ( .A0(weight_1[310]), .A1(n17787), .B0(weight_1[190]), .B1(
        n17790), .Y(n16761) );
  NAND4XL U20786 ( .A(n16764), .B(n16763), .C(n16762), .D(n16761), .Y(n16765)
         );
  NOR4XL U20787 ( .A(n16768), .B(n16767), .C(n16766), .D(n16765), .Y(n16769)
         );
  NAND2XL U20788 ( .A(n16770), .B(n16769), .Y(n16771) );
  OAI32XL U20789 ( .A0(n19182), .A1(n16773), .A2(n16772), .B0(cursor[6]), .B1(
        n16771), .Y(n16774) );
  NAND4XL U20790 ( .A(n16777), .B(n16776), .C(n16775), .D(n16774), .Y(n17162)
         );
  NAND2XL U20791 ( .A(n20645), .B(n17162), .Y(n17160) );
  NAND2BXL U20792 ( .AN(affine_1[24]), .B(n17160), .Y(
        DP_OP_5166J1_122_9881_n39) );
  AOI22XL U20793 ( .A0(n16734), .A1(weight_1[405]), .B0(n19097), .B1(
        weight_1[435]), .Y(n16781) );
  AOI22XL U20794 ( .A0(n21887), .A1(weight_1[417]), .B0(n19099), .B1(
        weight_1[429]), .Y(n16780) );
  AOI22XL U20795 ( .A0(n19098), .A1(weight_1[441]), .B0(n21954), .B1(
        weight_1[399]), .Y(n16779) );
  AOI22XL U20796 ( .A0(n22021), .A1(weight_1[411]), .B0(n19475), .B1(
        weight_1[423]), .Y(n16778) );
  NAND4XL U20797 ( .A(n16781), .B(n16780), .C(n16779), .D(n16778), .Y(n16784)
         );
  INVXL U20798 ( .A(weight_1[459]), .Y(n32478) );
  INVXL U20799 ( .A(weight_1[447]), .Y(n32484) );
  OAI22XL U20800 ( .A0(n32478), .A1(n17837), .B0(n32484), .B1(n17690), .Y(
        n16783) );
  INVXL U20801 ( .A(weight_1[465]), .Y(n32473) );
  INVXL U20802 ( .A(weight_1[453]), .Y(n32483) );
  OAI22XL U20803 ( .A0(n32473), .A1(n17747), .B0(n32483), .B1(n17746), .Y(
        n16782) );
  AOI211XL U20804 ( .A0(n17166), .A1(n16784), .B0(n16783), .C0(n16782), .Y(
        n16833) );
  INVXL U20805 ( .A(weight_1[471]), .Y(n32461) );
  INVXL U20806 ( .A(weight_1[9]), .Y(n32401) );
  INVXL U20807 ( .A(n17444), .Y(n17248) );
  OAI22XL U20808 ( .A0(n32461), .A1(n17846), .B0(n32401), .B1(n17248), .Y(
        n16831) );
  AOI22XL U20809 ( .A0(weight_1[309]), .A1(n17787), .B0(weight_1[147]), .B1(
        n17875), .Y(n16788) );
  AOI22XL U20810 ( .A0(weight_1[285]), .A1(n17802), .B0(weight_1[27]), .B1(
        n17893), .Y(n16787) );
  AOI22XL U20811 ( .A0(n21766), .A1(weight_1[321]), .B0(weight_1[249]), .B1(
        n17797), .Y(n16786) );
  AOI22XL U20812 ( .A0(weight_1[279]), .A1(n17877), .B0(weight_1[117]), .B1(
        n17876), .Y(n16785) );
  NAND4XL U20813 ( .A(n16788), .B(n16787), .C(n16786), .D(n16785), .Y(n16804)
         );
  AOI22XL U20814 ( .A0(weight_1[51]), .A1(n17803), .B0(weight_1[33]), .B1(
        n17873), .Y(n16792) );
  AOI22XL U20815 ( .A0(weight_1[135]), .A1(n17895), .B0(weight_1[69]), .B1(
        n17883), .Y(n16791) );
  AOI22XL U20816 ( .A0(weight_1[129]), .A1(n17801), .B0(weight_1[105]), .B1(
        n17885), .Y(n16790) );
  AOI22XL U20817 ( .A0(weight_1[189]), .A1(n17790), .B0(weight_1[75]), .B1(
        n17865), .Y(n16789) );
  NAND4XL U20818 ( .A(n16792), .B(n16791), .C(n16790), .D(n16789), .Y(n16803)
         );
  AOI22XL U20819 ( .A0(weight_1[387]), .A1(n17821), .B0(weight_1[297]), .B1(
        n17826), .Y(n16796) );
  AOI22XL U20820 ( .A0(weight_1[369]), .A1(n17825), .B0(weight_1[351]), .B1(
        n17812), .Y(n16795) );
  AOI22XL U20821 ( .A0(weight_1[345]), .A1(n17823), .B0(weight_1[201]), .B1(
        n17813), .Y(n16794) );
  AOI22XL U20822 ( .A0(weight_1[339]), .A1(n17814), .B0(weight_1[153]), .B1(
        n17822), .Y(n16793) );
  NAND4XL U20823 ( .A(n16796), .B(n16795), .C(n16794), .D(n16793), .Y(n16802)
         );
  AOI22XL U20824 ( .A0(weight_1[381]), .A1(n17810), .B0(weight_1[159]), .B1(
        n17868), .Y(n16800) );
  AOI22XL U20825 ( .A0(weight_1[375]), .A1(n17809), .B0(weight_1[363]), .B1(
        n17827), .Y(n16799) );
  AOI22XL U20826 ( .A0(weight_1[357]), .A1(n17816), .B0(weight_1[243]), .B1(
        n17815), .Y(n16798) );
  AOI22XL U20827 ( .A0(weight_1[237]), .A1(n17824), .B0(weight_1[231]), .B1(
        n17811), .Y(n16797) );
  NAND4XL U20828 ( .A(n16800), .B(n16799), .C(n16798), .D(n16797), .Y(n16801)
         );
  NOR4XL U20829 ( .A(n16804), .B(n16803), .C(n16802), .D(n16801), .Y(n16829)
         );
  AOI22XL U20830 ( .A0(weight_1[393]), .A1(n17800), .B0(weight_1[267]), .B1(
        n17788), .Y(n16808) );
  AOI22XL U20831 ( .A0(weight_1[171]), .A1(n17888), .B0(weight_1[99]), .B1(
        n17897), .Y(n16807) );
  AOI22XL U20832 ( .A0(weight_1[225]), .A1(n17878), .B0(weight_1[177]), .B1(
        n17899), .Y(n16806) );
  AOI22XL U20833 ( .A0(n16744), .A1(weight_1[87]), .B0(weight_1[45]), .B1(
        n17874), .Y(n16805) );
  NAND4XL U20834 ( .A(n16808), .B(n16807), .C(n16806), .D(n16805), .Y(n16824)
         );
  AOI22XL U20835 ( .A0(weight_1[261]), .A1(n17886), .B0(weight_1[81]), .B1(
        n17799), .Y(n16812) );
  AOI22XL U20836 ( .A0(weight_1[207]), .A1(n17884), .B0(weight_1[195]), .B1(
        n17866), .Y(n16811) );
  AOI22XL U20837 ( .A0(weight_1[255]), .A1(n17896), .B0(weight_1[213]), .B1(
        n17898), .Y(n16810) );
  AOI22XL U20838 ( .A0(weight_1[63]), .A1(n17791), .B0(weight_1[57]), .B1(
        n17789), .Y(n16809) );
  NAND4XL U20839 ( .A(n16812), .B(n16811), .C(n16810), .D(n16809), .Y(n16823)
         );
  AOI22XL U20840 ( .A0(weight_1[291]), .A1(n17900), .B0(weight_1[273]), .B1(
        n17864), .Y(n16816) );
  AOI22XL U20841 ( .A0(n21764), .A1(weight_1[21]), .B0(n21748), .B1(
        weight_1[315]), .Y(n16815) );
  AOI22XL U20842 ( .A0(n26082), .A1(weight_1[327]), .B0(n21999), .B1(
        weight_1[93]), .Y(n16814) );
  AOI22XL U20843 ( .A0(n26059), .A1(weight_1[333]), .B0(weight_1[123]), .B1(
        n17792), .Y(n16813) );
  NAND4XL U20844 ( .A(n16816), .B(n16815), .C(n16814), .D(n16813), .Y(n16822)
         );
  AOI22XL U20845 ( .A0(weight_1[303]), .A1(n17798), .B0(weight_1[39]), .B1(
        n17867), .Y(n16820) );
  AOI22XL U20846 ( .A0(weight_1[183]), .A1(n16724), .B0(weight_1[141]), .B1(
        n17894), .Y(n16819) );
  AOI22XL U20847 ( .A0(n21762), .A1(weight_1[15]), .B0(weight_1[111]), .B1(
        n17887), .Y(n16818) );
  AOI22XL U20848 ( .A0(weight_1[219]), .A1(n17804), .B0(weight_1[165]), .B1(
        n17863), .Y(n16817) );
  NAND4XL U20849 ( .A(n16820), .B(n16819), .C(n16818), .D(n16817), .Y(n16821)
         );
  NOR4XL U20850 ( .A(n16824), .B(n16823), .C(n16822), .D(n16821), .Y(n16828)
         );
  INVXL U20851 ( .A(weight_1[195]), .Y(n32729) );
  INVXL U20852 ( .A(weight_1[477]), .Y(n32464) );
  INVXL U20853 ( .A(weight_1[393]), .Y(n32501) );
  OAI22XL U20854 ( .A0(n21536), .A1(n32464), .B0(n32501), .B1(n17391), .Y(
        n16825) );
  AOI211XL U20855 ( .A0(n17821), .A1(weight_1[3]), .B0(n16826), .C0(n16825), 
        .Y(n16827) );
  AOI32XL U20856 ( .A0(n16829), .A1(n19182), .A2(n16828), .B0(cursor[6]), .B1(
        n16827), .Y(n16830) );
  AOI211XL U20857 ( .A0(weight_1[483]), .A1(n17068), .B0(n16831), .C0(n16830), 
        .Y(n16832) );
  NAND2XL U20858 ( .A(n16833), .B(n16832), .Y(n17161) );
  AOI22XL U20859 ( .A0(counter[1]), .A1(pool[133]), .B0(counter[0]), .B1(
        pool[128]), .Y(n16854) );
  AOI22XL U20860 ( .A0(pool[53]), .A1(n17011), .B0(pool[43]), .B1(n17010), .Y(
        n16853) );
  INVXL U20861 ( .A(pool[58]), .Y(n24687) );
  INVXL U20862 ( .A(n16676), .Y(n17025) );
  INVXL U20863 ( .A(pool[73]), .Y(n26351) );
  OAI22XL U20864 ( .A0(n19227), .A1(n24687), .B0(n17025), .B1(n26351), .Y(
        n16835) );
  INVXL U20865 ( .A(pool[78]), .Y(n27370) );
  INVXL U20866 ( .A(pool[68]), .Y(n22050) );
  OAI22XL U20867 ( .A0(n18172), .A1(n27370), .B0(n18174), .B1(n22050), .Y(
        n16834) );
  INVXL U20868 ( .A(n18159), .Y(n17014) );
  INVXL U20869 ( .A(pool[48]), .Y(n25445) );
  OAI22XL U20870 ( .A0(n16836), .A1(n19247), .B0(n17014), .B1(n25445), .Y(
        n16851) );
  INVXL U20871 ( .A(pool[13]), .Y(n28619) );
  INVXL U20872 ( .A(pool[3]), .Y(n25684) );
  OAI22XL U20873 ( .A0(n17028), .A1(n28619), .B0(n17027), .B1(n25684), .Y(
        n16840) );
  INVXL U20874 ( .A(pool[18]), .Y(n27977) );
  INVXL U20875 ( .A(pool[33]), .Y(n22797) );
  OAI22XL U20876 ( .A0(n19227), .A1(n27977), .B0(n17025), .B1(n22797), .Y(
        n16839) );
  INVXL U20877 ( .A(pool[8]), .Y(n20159) );
  INVXL U20878 ( .A(pool[23]), .Y(n22097) );
  OAI22XL U20879 ( .A0(n17029), .A1(n20159), .B0(n17026), .B1(n22097), .Y(
        n16838) );
  INVXL U20880 ( .A(pool[38]), .Y(n20612) );
  INVXL U20881 ( .A(pool[28]), .Y(n30645) );
  OAI22XL U20882 ( .A0(n18172), .A1(n20612), .B0(n18174), .B1(n30645), .Y(
        n16837) );
  NOR4XL U20883 ( .A(n16840), .B(n16839), .C(n16838), .D(n16837), .Y(n16849)
         );
  OAI31XL U20884 ( .A0(pool[63]), .A1(pool[123]), .A2(pool[103]), .B0(n19228), 
        .Y(n16841) );
  NAND2XL U20885 ( .A(n16854), .B(n16841), .Y(n16847) );
  INVXL U20886 ( .A(n20605), .Y(n17018) );
  INVXL U20887 ( .A(pool[83]), .Y(n26119) );
  INVXL U20888 ( .A(pool[123]), .Y(n26705) );
  OAI22XL U20889 ( .A0(n17018), .A1(n26119), .B0(n26705), .B1(n17017), .Y(
        n16846) );
  AOI222XL U20890 ( .A0(n19006), .A1(pool[88]), .B0(n19007), .B1(pool[103]), 
        .C0(n19005), .C1(pool[93]), .Y(n16844) );
  AOI22XL U20891 ( .A0(n19008), .A1(pool[118]), .B0(n19004), .B1(pool[108]), 
        .Y(n16843) );
  AOI22XL U20892 ( .A0(n19009), .A1(pool[98]), .B0(n16676), .B1(pool[113]), 
        .Y(n16842) );
  OAI211XL U20893 ( .A0(counter[3]), .A1(n16844), .B0(n16843), .C0(n16842), 
        .Y(n16845) );
  AOI211XL U20894 ( .A0(n20363), .A1(n16847), .B0(n16846), .C0(n16845), .Y(
        n16848) );
  OAI22XL U20895 ( .A0(n16849), .A1(n18156), .B0(n16848), .B1(n20600), .Y(
        n16850) );
  AOI211XL U20896 ( .A0(pool[63]), .A1(n17038), .B0(n16851), .C0(n16850), .Y(
        n16852) );
  AOI22XL U20897 ( .A0(weight_1[218]), .A1(n17804), .B0(weight_1[68]), .B1(
        n17883), .Y(n16858) );
  AOI22XL U20898 ( .A0(weight_1[188]), .A1(n17790), .B0(weight_1[80]), .B1(
        n17799), .Y(n16857) );
  AOI22XL U20899 ( .A0(n21762), .A1(weight_1[14]), .B0(n21766), .B1(
        weight_1[320]), .Y(n16856) );
  AOI22XL U20900 ( .A0(weight_1[56]), .A1(n17789), .B0(weight_1[32]), .B1(
        n17873), .Y(n16855) );
  NAND4XL U20901 ( .A(n16858), .B(n16857), .C(n16856), .D(n16855), .Y(n16874)
         );
  AOI22XL U20902 ( .A0(weight_1[302]), .A1(n17798), .B0(weight_1[44]), .B1(
        n17874), .Y(n16862) );
  AOI22XL U20903 ( .A0(weight_1[284]), .A1(n17802), .B0(weight_1[158]), .B1(
        n17868), .Y(n16861) );
  AOI22XL U20904 ( .A0(weight_1[260]), .A1(n17886), .B0(weight_1[182]), .B1(
        n16724), .Y(n16860) );
  AOI22XL U20905 ( .A0(n21999), .A1(weight_1[92]), .B0(weight_1[272]), .B1(
        n17864), .Y(n16859) );
  NAND4XL U20906 ( .A(n16862), .B(n16861), .C(n16860), .D(n16859), .Y(n16873)
         );
  AOI22XL U20907 ( .A0(weight_1[368]), .A1(n17825), .B0(weight_1[242]), .B1(
        n17815), .Y(n16866) );
  AOI22XL U20908 ( .A0(weight_1[362]), .A1(n17827), .B0(weight_1[200]), .B1(
        n17813), .Y(n16865) );
  AOI22XL U20909 ( .A0(weight_1[386]), .A1(n17821), .B0(weight_1[236]), .B1(
        n17824), .Y(n16864) );
  AOI22XL U20910 ( .A0(weight_1[230]), .A1(n17811), .B0(weight_1[152]), .B1(
        n17822), .Y(n16863) );
  NAND4XL U20911 ( .A(n16866), .B(n16865), .C(n16864), .D(n16863), .Y(n16872)
         );
  AOI22XL U20912 ( .A0(weight_1[350]), .A1(n17812), .B0(weight_1[290]), .B1(
        n17900), .Y(n16870) );
  AOI22XL U20913 ( .A0(weight_1[338]), .A1(n17814), .B0(weight_1[296]), .B1(
        n17826), .Y(n16869) );
  AOI22XL U20914 ( .A0(weight_1[356]), .A1(n17816), .B0(weight_1[344]), .B1(
        n17823), .Y(n16868) );
  AOI22XL U20915 ( .A0(weight_1[380]), .A1(n17810), .B0(weight_1[374]), .B1(
        n17809), .Y(n16867) );
  NAND4XL U20916 ( .A(n16870), .B(n16869), .C(n16868), .D(n16867), .Y(n16871)
         );
  NOR4XL U20917 ( .A(n16874), .B(n16873), .C(n16872), .D(n16871), .Y(n16909)
         );
  INVXL U20918 ( .A(weight_1[476]), .Y(n32679) );
  INVXL U20919 ( .A(weight_1[8]), .Y(n32378) );
  OAI22XL U20920 ( .A0(n32679), .A1(n17694), .B0(n32378), .B1(n17248), .Y(
        n16886) );
  INVXL U20921 ( .A(n17746), .Y(n17849) );
  AOI22XL U20922 ( .A0(weight_1[470]), .A1(n17691), .B0(weight_1[452]), .B1(
        n17849), .Y(n16884) );
  INVXL U20923 ( .A(weight_1[194]), .Y(n32743) );
  INVXL U20924 ( .A(weight_1[2]), .Y(n32371) );
  OAI22XL U20925 ( .A0(n32743), .A1(n17143), .B0(n32371), .B1(n17188), .Y(
        n16875) );
  AOI22XL U20926 ( .A0(cursor[6]), .A1(n16875), .B0(weight_1[464]), .B1(n17852), .Y(n16883) );
  AOI22XL U20927 ( .A0(n19097), .A1(weight_1[434]), .B0(n19099), .B1(
        weight_1[428]), .Y(n16879) );
  AOI22XL U20928 ( .A0(n16734), .A1(weight_1[404]), .B0(n21954), .B1(
        weight_1[398]), .Y(n16878) );
  AOI22XL U20929 ( .A0(n19098), .A1(weight_1[440]), .B0(n19475), .B1(
        weight_1[422]), .Y(n16877) );
  AOI22XL U20930 ( .A0(n22021), .A1(weight_1[410]), .B0(n21887), .B1(
        weight_1[416]), .Y(n16876) );
  NAND4XL U20931 ( .A(n16879), .B(n16878), .C(n16877), .D(n16876), .Y(n16880)
         );
  AOI22XL U20932 ( .A0(weight_1[458]), .A1(n17753), .B0(n17166), .B1(n16880), 
        .Y(n16882) );
  AOI22XL U20933 ( .A0(weight_1[446]), .A1(n17848), .B0(weight_1[392]), .B1(
        n17454), .Y(n16881) );
  NAND4XL U20934 ( .A(n16884), .B(n16883), .C(n16882), .D(n16881), .Y(n16885)
         );
  AOI211XL U20935 ( .A0(weight_1[482]), .A1(n17068), .B0(n16886), .C0(n16885), 
        .Y(n16908) );
  AOI22XL U20936 ( .A0(weight_1[140]), .A1(n17894), .B0(weight_1[50]), .B1(
        n17803), .Y(n16890) );
  AOI22XL U20937 ( .A0(weight_1[98]), .A1(n17897), .B0(weight_1[74]), .B1(
        n17865), .Y(n16889) );
  AOI22XL U20938 ( .A0(weight_1[392]), .A1(n17800), .B0(weight_1[104]), .B1(
        n17885), .Y(n16888) );
  AOI22XL U20939 ( .A0(weight_1[254]), .A1(n17896), .B0(weight_1[110]), .B1(
        n17887), .Y(n16887) );
  NAND4XL U20940 ( .A(n16890), .B(n16889), .C(n16888), .D(n16887), .Y(n16906)
         );
  AOI22XL U20941 ( .A0(weight_1[266]), .A1(n17788), .B0(weight_1[116]), .B1(
        n17876), .Y(n16894) );
  AOI22XL U20942 ( .A0(weight_1[194]), .A1(n17866), .B0(weight_1[128]), .B1(
        n17801), .Y(n16893) );
  AOI22XL U20943 ( .A0(weight_1[248]), .A1(n17797), .B0(weight_1[170]), .B1(
        n17888), .Y(n16892) );
  AOI22XL U20944 ( .A0(weight_1[224]), .A1(n17878), .B0(weight_1[38]), .B1(
        n17867), .Y(n16891) );
  NAND4XL U20945 ( .A(n16894), .B(n16893), .C(n16892), .D(n16891), .Y(n16905)
         );
  AOI22XL U20946 ( .A0(weight_1[308]), .A1(n17787), .B0(weight_1[146]), .B1(
        n17875), .Y(n16898) );
  AOI22XL U20947 ( .A0(n26082), .A1(weight_1[326]), .B0(weight_1[134]), .B1(
        n17895), .Y(n16897) );
  AOI22XL U20948 ( .A0(n26059), .A1(weight_1[332]), .B0(weight_1[62]), .B1(
        n17791), .Y(n16896) );
  AOI22XL U20949 ( .A0(weight_1[212]), .A1(n17898), .B0(weight_1[176]), .B1(
        n17899), .Y(n16895) );
  NAND4XL U20950 ( .A(n16898), .B(n16897), .C(n16896), .D(n16895), .Y(n16904)
         );
  AOI22XL U20951 ( .A0(n21764), .A1(weight_1[20]), .B0(weight_1[26]), .B1(
        n17893), .Y(n16902) );
  AOI22XL U20952 ( .A0(n16744), .A1(weight_1[86]), .B0(weight_1[206]), .B1(
        n17884), .Y(n16901) );
  AOI22XL U20953 ( .A0(weight_1[164]), .A1(n17863), .B0(weight_1[122]), .B1(
        n17792), .Y(n16900) );
  AOI22XL U20954 ( .A0(n21748), .A1(weight_1[314]), .B0(weight_1[278]), .B1(
        n17877), .Y(n16899) );
  NAND4XL U20955 ( .A(n16902), .B(n16901), .C(n16900), .D(n16899), .Y(n16903)
         );
  NOR4XL U20956 ( .A(n16906), .B(n16905), .C(n16904), .D(n16903), .Y(n16907)
         );
  AOI32XL U20957 ( .A0(n16909), .A1(n16908), .A2(n16907), .B0(cursor[6]), .B1(
        n16908), .Y(n20613) );
  AND2XL U20958 ( .A(n20613), .B(n17918), .Y(DP_OP_5166J1_122_9881_n61) );
  INVXL U20959 ( .A(weight_1[468]), .Y(n26907) );
  AOI22XL U20960 ( .A0(weight_1[480]), .A1(n17068), .B0(weight_1[474]), .B1(
        n17842), .Y(n16965) );
  INVXL U20961 ( .A(weight_1[450]), .Y(n26867) );
  AOI22XL U20962 ( .A0(weight_1[456]), .A1(n17753), .B0(weight_1[444]), .B1(
        n17848), .Y(n16910) );
  OAI21XL U20963 ( .A0(n26867), .A1(n17746), .B0(n16910), .Y(n16963) );
  AOI22XL U20964 ( .A0(weight_1[282]), .A1(n17802), .B0(weight_1[108]), .B1(
        n17887), .Y(n16914) );
  AOI22XL U20965 ( .A0(weight_1[210]), .A1(n17898), .B0(weight_1[102]), .B1(
        n17885), .Y(n16913) );
  AOI22XL U20966 ( .A0(weight_1[288]), .A1(n17900), .B0(weight_1[66]), .B1(
        n17883), .Y(n16912) );
  AOI22XL U20967 ( .A0(n21762), .A1(weight_1[12]), .B0(weight_1[264]), .B1(
        n17788), .Y(n16911) );
  NAND4XL U20968 ( .A(n16914), .B(n16913), .C(n16912), .D(n16911), .Y(n16930)
         );
  AOI22XL U20969 ( .A0(n21999), .A1(weight_1[90]), .B0(weight_1[132]), .B1(
        n17895), .Y(n16918) );
  AOI22XL U20970 ( .A0(weight_1[258]), .A1(n17886), .B0(weight_1[174]), .B1(
        n17899), .Y(n16917) );
  AOI22XL U20971 ( .A0(weight_1[270]), .A1(n17864), .B0(weight_1[36]), .B1(
        n17867), .Y(n16916) );
  AOI22XL U20972 ( .A0(weight_1[186]), .A1(n17790), .B0(weight_1[156]), .B1(
        n17868), .Y(n16915) );
  NAND4XL U20973 ( .A(n16918), .B(n16917), .C(n16916), .D(n16915), .Y(n16929)
         );
  AOI22XL U20974 ( .A0(weight_1[366]), .A1(n17825), .B0(weight_1[354]), .B1(
        n17816), .Y(n16922) );
  AOI22XL U20975 ( .A0(weight_1[336]), .A1(n17814), .B0(weight_1[234]), .B1(
        n17824), .Y(n16921) );
  AOI22XL U20976 ( .A0(weight_1[348]), .A1(n17812), .B0(weight_1[228]), .B1(
        n17811), .Y(n16920) );
  AOI22XL U20977 ( .A0(weight_1[360]), .A1(n17827), .B0(weight_1[198]), .B1(
        n17813), .Y(n16919) );
  NAND4XL U20978 ( .A(n16922), .B(n16921), .C(n16920), .D(n16919), .Y(n16928)
         );
  AOI22XL U20979 ( .A0(weight_1[372]), .A1(n17809), .B0(weight_1[216]), .B1(
        n17804), .Y(n16926) );
  AOI22XL U20980 ( .A0(weight_1[294]), .A1(n17826), .B0(weight_1[150]), .B1(
        n17822), .Y(n16925) );
  AOI22XL U20981 ( .A0(weight_1[384]), .A1(n17821), .B0(weight_1[378]), .B1(
        n17810), .Y(n16924) );
  AOI22XL U20982 ( .A0(weight_1[342]), .A1(n17823), .B0(weight_1[240]), .B1(
        n17815), .Y(n16923) );
  NAND4XL U20983 ( .A(n16926), .B(n16925), .C(n16924), .D(n16923), .Y(n16927)
         );
  NOR4XL U20984 ( .A(n16930), .B(n16929), .C(n16928), .D(n16927), .Y(n16961)
         );
  AOI22XL U20985 ( .A0(weight_1[390]), .A1(n17800), .B0(weight_1[204]), .B1(
        n17884), .Y(n16934) );
  AOI22XL U20986 ( .A0(weight_1[276]), .A1(n17877), .B0(weight_1[42]), .B1(
        n17874), .Y(n16933) );
  AOI22XL U20987 ( .A0(n21748), .A1(weight_1[312]), .B0(weight_1[48]), .B1(
        n17803), .Y(n16932) );
  AOI22XL U20988 ( .A0(weight_1[252]), .A1(n17896), .B0(weight_1[96]), .B1(
        n17897), .Y(n16931) );
  NAND4XL U20989 ( .A(n16934), .B(n16933), .C(n16932), .D(n16931), .Y(n16950)
         );
  AOI22XL U20990 ( .A0(n21764), .A1(weight_1[18]), .B0(weight_1[246]), .B1(
        n17797), .Y(n16938) );
  AOI22XL U20991 ( .A0(weight_1[192]), .A1(n17866), .B0(weight_1[54]), .B1(
        n17789), .Y(n16937) );
  AOI22XL U20992 ( .A0(weight_1[120]), .A1(n17792), .B0(weight_1[78]), .B1(
        n17799), .Y(n16936) );
  AOI22XL U20993 ( .A0(weight_1[162]), .A1(n17863), .B0(weight_1[144]), .B1(
        n17875), .Y(n16935) );
  NAND4XL U20994 ( .A(n16938), .B(n16937), .C(n16936), .D(n16935), .Y(n16949)
         );
  AOI22XL U20995 ( .A0(weight_1[168]), .A1(n17888), .B0(weight_1[138]), .B1(
        n17894), .Y(n16942) );
  AOI22XL U20996 ( .A0(n21766), .A1(weight_1[318]), .B0(weight_1[72]), .B1(
        n17865), .Y(n16941) );
  AOI22XL U20997 ( .A0(weight_1[30]), .A1(n17873), .B0(weight_1[24]), .B1(
        n17893), .Y(n16940) );
  AOI22XL U20998 ( .A0(weight_1[126]), .A1(n17801), .B0(weight_1[114]), .B1(
        n17876), .Y(n16939) );
  NAND4XL U20999 ( .A(n16942), .B(n16941), .C(n16940), .D(n16939), .Y(n16948)
         );
  AOI22XL U21000 ( .A0(n16744), .A1(weight_1[84]), .B0(weight_1[222]), .B1(
        n17878), .Y(n16946) );
  AOI22XL U21001 ( .A0(weight_1[300]), .A1(n17798), .B0(weight_1[180]), .B1(
        n16724), .Y(n16945) );
  AOI22XL U21002 ( .A0(n26059), .A1(weight_1[330]), .B0(weight_1[306]), .B1(
        n17787), .Y(n16944) );
  AOI22XL U21003 ( .A0(n26082), .A1(weight_1[324]), .B0(weight_1[60]), .B1(
        n17791), .Y(n16943) );
  NAND4XL U21004 ( .A(n16946), .B(n16945), .C(n16944), .D(n16943), .Y(n16947)
         );
  NOR4XL U21005 ( .A(n16950), .B(n16949), .C(n16948), .D(n16947), .Y(n16960)
         );
  INVXL U21006 ( .A(weight_1[192]), .Y(n26868) );
  INVXL U21007 ( .A(weight_1[6]), .Y(n32724) );
  OAI22XL U21008 ( .A0(n26868), .A1(n17143), .B0(n32724), .B1(n16951), .Y(
        n16958) );
  INVXL U21009 ( .A(weight_1[414]), .Y(n26891) );
  INVXL U21010 ( .A(weight_1[426]), .Y(n26871) );
  OAI22XL U21011 ( .A0(n21810), .A1(n26891), .B0(n17173), .B1(n26871), .Y(
        n16955) );
  INVXL U21012 ( .A(weight_1[402]), .Y(n26911) );
  INVXL U21013 ( .A(weight_1[438]), .Y(n26885) );
  OAI22XL U21014 ( .A0(n21944), .A1(n26911), .B0(n17170), .B1(n26885), .Y(
        n16954) );
  INVXL U21015 ( .A(weight_1[420]), .Y(n26857) );
  INVXL U21016 ( .A(weight_1[396]), .Y(n26912) );
  OAI22XL U21017 ( .A0(n17165), .A1(n26857), .B0(n16669), .B1(n26912), .Y(
        n16953) );
  INVXL U21018 ( .A(weight_1[408]), .Y(n26892) );
  INVXL U21019 ( .A(weight_1[432]), .Y(n26886) );
  OAI22XL U21020 ( .A0(n19416), .A1(n26892), .B0(n20726), .B1(n26886), .Y(
        n16952) );
  NOR4XL U21021 ( .A(n16955), .B(n16954), .C(n16953), .D(n16952), .Y(n16956)
         );
  INVXL U21022 ( .A(weight_1[0]), .Y(n32414) );
  OAI22XL U21023 ( .A0(n16956), .A1(n35159), .B0(n32414), .B1(n17188), .Y(
        n16957) );
  AOI211XL U21024 ( .A0(weight_1[390]), .A1(n17813), .B0(n16958), .C0(n16957), 
        .Y(n16959) );
  AOI32XL U21025 ( .A0(n16961), .A1(n19182), .A2(n16960), .B0(cursor[6]), .B1(
        n16959), .Y(n16962) );
  AOI211XL U21026 ( .A0(weight_1[462]), .A1(n17852), .B0(n16963), .C0(n16962), 
        .Y(n16964) );
  OAI211XL U21027 ( .A0(n26907), .A1(n17846), .B0(n16965), .C0(n16964), .Y(
        n20624) );
  AND2XL U21028 ( .A(n20624), .B(n17918), .Y(DP_OP_5166J1_122_9881_n63) );
  AOI22XL U21029 ( .A0(counter[1]), .A1(pool[132]), .B0(counter[0]), .B1(
        pool[127]), .Y(n16986) );
  AOI22XL U21030 ( .A0(pool[52]), .A1(n17011), .B0(pool[42]), .B1(n17010), .Y(
        n16985) );
  INVXL U21031 ( .A(pool[67]), .Y(n34891) );
  INVXL U21032 ( .A(pool[57]), .Y(n34877) );
  INVXL U21033 ( .A(pool[77]), .Y(n34900) );
  OAI22XL U21034 ( .A0(n19227), .A1(n34877), .B0(n18172), .B1(n34900), .Y(
        n16966) );
  AOI211XL U21035 ( .A0(pool[72]), .A1(n16676), .B0(n16967), .C0(n16966), .Y(
        n16968) );
  INVXL U21036 ( .A(pool[47]), .Y(n34867) );
  OAI22XL U21037 ( .A0(n16968), .A1(n19247), .B0(n17014), .B1(n34867), .Y(
        n16983) );
  INVXL U21038 ( .A(pool[7]), .Y(n34801) );
  INVXL U21039 ( .A(pool[27]), .Y(n34820) );
  OAI22XL U21040 ( .A0(n17029), .A1(n34801), .B0(n18174), .B1(n34820), .Y(
        n16972) );
  INVXL U21041 ( .A(pool[17]), .Y(n34811) );
  INVXL U21042 ( .A(pool[2]), .Y(n34793) );
  OAI22XL U21043 ( .A0(n19227), .A1(n34811), .B0(n17027), .B1(n34793), .Y(
        n16971) );
  INVXL U21044 ( .A(pool[37]), .Y(n34843) );
  INVXL U21045 ( .A(pool[32]), .Y(n34838) );
  OAI22XL U21046 ( .A0(n18172), .A1(n34843), .B0(n17025), .B1(n34838), .Y(
        n16970) );
  INVXL U21047 ( .A(pool[22]), .Y(n34816) );
  INVXL U21048 ( .A(pool[12]), .Y(n34805) );
  OAI22XL U21049 ( .A0(n17026), .A1(n34816), .B0(n17028), .B1(n34805), .Y(
        n16969) );
  NOR4XL U21050 ( .A(n16972), .B(n16971), .C(n16970), .D(n16969), .Y(n16981)
         );
  OAI31XL U21051 ( .A0(pool[62]), .A1(pool[122]), .A2(pool[102]), .B0(n19228), 
        .Y(n16973) );
  NAND2XL U21052 ( .A(n16986), .B(n16973), .Y(n16979) );
  INVXL U21053 ( .A(pool[82]), .Y(n34925) );
  INVXL U21054 ( .A(pool[122]), .Y(n35021) );
  OAI22XL U21055 ( .A0(n17018), .A1(n34925), .B0(n35021), .B1(n17017), .Y(
        n16978) );
  AOI222XL U21056 ( .A0(n19006), .A1(pool[87]), .B0(n19007), .B1(pool[102]), 
        .C0(n19005), .C1(pool[92]), .Y(n16976) );
  AOI22XL U21057 ( .A0(n19009), .A1(pool[97]), .B0(n19008), .B1(pool[117]), 
        .Y(n16975) );
  AOI22XL U21058 ( .A0(n19004), .A1(pool[107]), .B0(n16676), .B1(pool[112]), 
        .Y(n16974) );
  OAI211XL U21059 ( .A0(counter[3]), .A1(n16976), .B0(n16975), .C0(n16974), 
        .Y(n16977) );
  AOI211XL U21060 ( .A0(n20363), .A1(n16979), .B0(n16978), .C0(n16977), .Y(
        n16980) );
  OAI22XL U21061 ( .A0(n16981), .A1(n18156), .B0(n16980), .B1(n20600), .Y(
        n16982) );
  AOI211XL U21062 ( .A0(pool[62]), .A1(n17038), .B0(n16983), .C0(n16982), .Y(
        n16984) );
  AND2XL U21063 ( .A(n17162), .B(n20646), .Y(DP_OP_5166J1_122_9881_n65) );
  AND2XL U21064 ( .A(n17161), .B(n20646), .Y(DP_OP_5166J1_122_9881_n66) );
  AND2XL U21065 ( .A(n20613), .B(n20646), .Y(DP_OP_5166J1_122_9881_n67) );
  AOI22XL U21066 ( .A0(counter[1]), .A1(pool[131]), .B0(counter[0]), .B1(
        pool[126]), .Y(n17009) );
  AOI22XL U21067 ( .A0(pool[51]), .A1(n17011), .B0(pool[41]), .B1(n17010), .Y(
        n17008) );
  AOI22XL U21068 ( .A0(n19008), .A1(pool[36]), .B0(n19005), .B1(pool[11]), .Y(
        n16991) );
  AOI22XL U21069 ( .A0(n19007), .A1(pool[21]), .B0(n16987), .B1(pool[1]), .Y(
        n16990) );
  AOI22XL U21070 ( .A0(n19009), .A1(pool[16]), .B0(n16676), .B1(pool[31]), .Y(
        n16989) );
  AOI22XL U21071 ( .A0(n19006), .A1(pool[6]), .B0(n19004), .B1(pool[26]), .Y(
        n16988) );
  NAND4XL U21072 ( .A(n16991), .B(n16990), .C(n16989), .D(n16988), .Y(n17005)
         );
  AOI22XL U21073 ( .A0(n19009), .A1(pool[96]), .B0(n16676), .B1(pool[111]), 
        .Y(n16999) );
  OAI31XL U21074 ( .A0(pool[61]), .A1(pool[121]), .A2(pool[101]), .B0(n19228), 
        .Y(n16992) );
  AOI21XL U21075 ( .A0(n17009), .A1(n16992), .B0(n18170), .Y(n16994) );
  INVXL U21076 ( .A(pool[106]), .Y(n35005) );
  INVXL U21077 ( .A(pool[121]), .Y(n26703) );
  OAI22XL U21078 ( .A0(n18174), .A1(n35005), .B0(n26703), .B1(n17017), .Y(
        n16993) );
  AOI211XL U21079 ( .A0(pool[116]), .A1(n19008), .B0(n16994), .C0(n16993), .Y(
        n16998) );
  INVXL U21080 ( .A(pool[101]), .Y(n34996) );
  INVXL U21081 ( .A(pool[81]), .Y(n26114) );
  OAI22XL U21082 ( .A0(n17026), .A1(n34996), .B0(n17027), .B1(n26114), .Y(
        n16996) );
  INVXL U21083 ( .A(pool[86]), .Y(n22199) );
  INVXL U21084 ( .A(pool[91]), .Y(n27068) );
  OAI22XL U21085 ( .A0(n17029), .A1(n22199), .B0(n17028), .B1(n27068), .Y(
        n16995) );
  OAI21XL U21086 ( .A0(n16996), .A1(n16995), .B0(n19247), .Y(n16997) );
  AOI31XL U21087 ( .A0(n16999), .A1(n16998), .A2(n16997), .B0(n20600), .Y(
        n17004) );
  AOI22XL U21088 ( .A0(n19008), .A1(pool[76]), .B0(n19004), .B1(pool[66]), .Y(
        n17002) );
  AOI22XL U21089 ( .A0(n19009), .A1(pool[56]), .B0(n16676), .B1(pool[71]), .Y(
        n17001) );
  AOI22XL U21090 ( .A0(n18159), .A1(pool[46]), .B0(pool[61]), .B1(n17038), .Y(
        n17000) );
  AOI31XL U21091 ( .A0(n17002), .A1(n17001), .A2(n17000), .B0(n19247), .Y(
        n17003) );
  AOI211XL U21092 ( .A0(n17006), .A1(n17005), .B0(n17004), .C0(n17003), .Y(
        n17007) );
  AND2XL U21093 ( .A(n20613), .B(n20648), .Y(DP_OP_5166J1_122_9881_n73) );
  AOI22XL U21094 ( .A0(counter[1]), .A1(pool[134]), .B0(counter[0]), .B1(
        pool[129]), .Y(n17041) );
  AOI22XL U21095 ( .A0(pool[54]), .A1(n17011), .B0(pool[44]), .B1(n17010), .Y(
        n17040) );
  INVXL U21096 ( .A(pool[59]), .Y(n34879) );
  INVXL U21097 ( .A(pool[79]), .Y(n27372) );
  OAI22XL U21098 ( .A0(n19227), .A1(n34879), .B0(n18172), .B1(n27372), .Y(
        n17013) );
  INVXL U21099 ( .A(pool[69]), .Y(n22052) );
  INVXL U21100 ( .A(pool[74]), .Y(n26349) );
  OAI22XL U21101 ( .A0(n18174), .A1(n22052), .B0(n17025), .B1(n26349), .Y(
        n17012) );
  INVXL U21102 ( .A(pool[49]), .Y(n25443) );
  OAI22XL U21103 ( .A0(n17015), .A1(n19247), .B0(n17014), .B1(n25443), .Y(
        n17037) );
  OAI31XL U21104 ( .A0(pool[64]), .A1(pool[124]), .A2(pool[104]), .B0(n19228), 
        .Y(n17016) );
  NAND2XL U21105 ( .A(n17041), .B(n17016), .Y(n17024) );
  INVXL U21106 ( .A(pool[84]), .Y(n26116) );
  INVXL U21107 ( .A(pool[124]), .Y(n26708) );
  OAI22XL U21108 ( .A0(n17018), .A1(n26116), .B0(n26708), .B1(n17017), .Y(
        n17023) );
  AOI222XL U21109 ( .A0(n19006), .A1(pool[89]), .B0(n19007), .B1(pool[104]), 
        .C0(n19005), .C1(pool[94]), .Y(n17021) );
  AOI22XL U21110 ( .A0(n19009), .A1(pool[99]), .B0(n16676), .B1(pool[114]), 
        .Y(n17020) );
  AOI22XL U21111 ( .A0(n19008), .A1(pool[119]), .B0(n19004), .B1(pool[109]), 
        .Y(n17019) );
  OAI211XL U21112 ( .A0(counter[3]), .A1(n17021), .B0(n17020), .C0(n17019), 
        .Y(n17022) );
  AOI211XL U21113 ( .A0(n20363), .A1(n17024), .B0(n17023), .C0(n17022), .Y(
        n17035) );
  INVXL U21114 ( .A(pool[19]), .Y(n27979) );
  INVXL U21115 ( .A(pool[34]), .Y(n22799) );
  OAI22XL U21116 ( .A0(n19227), .A1(n27979), .B0(n17025), .B1(n22799), .Y(
        n17033) );
  INVXL U21117 ( .A(pool[29]), .Y(n30647) );
  INVXL U21118 ( .A(pool[24]), .Y(n22095) );
  OAI22XL U21119 ( .A0(n18174), .A1(n30647), .B0(n17026), .B1(n22095), .Y(
        n17032) );
  INVXL U21120 ( .A(pool[39]), .Y(n20610) );
  INVXL U21121 ( .A(pool[4]), .Y(n34796) );
  OAI22XL U21122 ( .A0(n18172), .A1(n20610), .B0(n17027), .B1(n34796), .Y(
        n17031) );
  INVXL U21123 ( .A(pool[9]), .Y(n20161) );
  INVXL U21124 ( .A(pool[14]), .Y(n28617) );
  OAI22XL U21125 ( .A0(n17029), .A1(n20161), .B0(n17028), .B1(n28617), .Y(
        n17030) );
  NOR4XL U21126 ( .A(n17033), .B(n17032), .C(n17031), .D(n17030), .Y(n17034)
         );
  OAI22XL U21127 ( .A0(n17035), .A1(n20600), .B0(n17034), .B1(n18156), .Y(
        n17036) );
  AOI211XL U21128 ( .A0(pool[64]), .A1(n17038), .B0(n17037), .C0(n17036), .Y(
        n17039) );
  NAND2XL U21129 ( .A(n33554), .B(n20624), .Y(DP_OP_5166J1_122_9881_n57) );
  AOI22XL U21130 ( .A0(weight_1[269]), .A1(n17788), .B0(weight_1[209]), .B1(
        n17884), .Y(n17045) );
  AOI22XL U21131 ( .A0(n26059), .A1(weight_1[335]), .B0(weight_1[293]), .B1(
        n17900), .Y(n17044) );
  AOI22XL U21132 ( .A0(weight_1[125]), .A1(n17792), .B0(weight_1[107]), .B1(
        n17885), .Y(n17043) );
  AOI22XL U21133 ( .A0(weight_1[101]), .A1(n17897), .B0(weight_1[59]), .B1(
        n17789), .Y(n17042) );
  NAND4XL U21134 ( .A(n17045), .B(n17044), .C(n17043), .D(n17042), .Y(n17061)
         );
  AOI22XL U21135 ( .A0(weight_1[287]), .A1(n17802), .B0(weight_1[47]), .B1(
        n17874), .Y(n17049) );
  AOI22XL U21136 ( .A0(n21999), .A1(weight_1[95]), .B0(n21764), .B1(
        weight_1[23]), .Y(n17048) );
  AOI22XL U21137 ( .A0(weight_1[275]), .A1(n17864), .B0(weight_1[185]), .B1(
        n16724), .Y(n17047) );
  AOI22XL U21138 ( .A0(n21762), .A1(weight_1[17]), .B0(weight_1[173]), .B1(
        n17888), .Y(n17046) );
  NAND4XL U21139 ( .A(n17049), .B(n17048), .C(n17047), .D(n17046), .Y(n17060)
         );
  AOI22XL U21140 ( .A0(weight_1[377]), .A1(n17809), .B0(weight_1[371]), .B1(
        n17825), .Y(n17053) );
  AOI22XL U21141 ( .A0(weight_1[353]), .A1(n17812), .B0(weight_1[347]), .B1(
        n17823), .Y(n17052) );
  AOI22XL U21142 ( .A0(weight_1[341]), .A1(n17814), .B0(weight_1[155]), .B1(
        n17822), .Y(n17051) );
  AOI22XL U21143 ( .A0(weight_1[383]), .A1(n17810), .B0(weight_1[245]), .B1(
        n17815), .Y(n17050) );
  NAND4XL U21144 ( .A(n17053), .B(n17052), .C(n17051), .D(n17050), .Y(n17059)
         );
  AOI22XL U21145 ( .A0(weight_1[299]), .A1(n17826), .B0(weight_1[119]), .B1(
        n17876), .Y(n17057) );
  AOI22XL U21146 ( .A0(weight_1[359]), .A1(n17816), .B0(weight_1[203]), .B1(
        n17813), .Y(n17056) );
  AOI22XL U21147 ( .A0(weight_1[389]), .A1(n17821), .B0(weight_1[239]), .B1(
        n17824), .Y(n17055) );
  AOI22XL U21148 ( .A0(weight_1[365]), .A1(n17827), .B0(weight_1[233]), .B1(
        n17811), .Y(n17054) );
  NAND4XL U21149 ( .A(n17057), .B(n17056), .C(n17055), .D(n17054), .Y(n17058)
         );
  NOR4XL U21150 ( .A(n17061), .B(n17060), .C(n17059), .D(n17058), .Y(n17098)
         );
  AOI22XL U21151 ( .A0(n19098), .A1(weight_1[443]), .B0(n19475), .B1(
        weight_1[425]), .Y(n17065) );
  AOI22XL U21152 ( .A0(n22021), .A1(weight_1[413]), .B0(n21954), .B1(
        weight_1[401]), .Y(n17064) );
  AOI22XL U21153 ( .A0(n19097), .A1(weight_1[437]), .B0(n19099), .B1(
        weight_1[431]), .Y(n17063) );
  AOI22XL U21154 ( .A0(n16734), .A1(weight_1[407]), .B0(n21887), .B1(
        weight_1[419]), .Y(n17062) );
  NAND4XL U21155 ( .A(n17065), .B(n17064), .C(n17063), .D(n17062), .Y(n17075)
         );
  AOI22XL U21156 ( .A0(weight_1[11]), .A1(n17800), .B0(weight_1[5]), .B1(
        n17821), .Y(n17067) );
  NAND2XL U21157 ( .A(weight_1[197]), .B(n17866), .Y(n17066) );
  AOI21XL U21158 ( .A0(n17067), .A1(n17066), .B0(n19182), .Y(n17074) );
  INVXL U21159 ( .A(weight_1[479]), .Y(n32930) );
  AOI22XL U21160 ( .A0(weight_1[485]), .A1(n17068), .B0(weight_1[395]), .B1(
        n17454), .Y(n17072) );
  INVXL U21161 ( .A(weight_1[455]), .Y(n32902) );
  INVXL U21162 ( .A(weight_1[449]), .Y(n32922) );
  OAI22XL U21163 ( .A0(n32902), .A1(n17746), .B0(n32922), .B1(n17690), .Y(
        n17070) );
  INVXL U21164 ( .A(weight_1[467]), .Y(n32906) );
  INVXL U21165 ( .A(weight_1[461]), .Y(n32901) );
  OAI22XL U21166 ( .A0(n32906), .A1(n17747), .B0(n32901), .B1(n17837), .Y(
        n17069) );
  AOI211XL U21167 ( .A0(weight_1[473]), .A1(n17691), .B0(n17070), .C0(n17069), 
        .Y(n17071) );
  OAI211XL U21168 ( .A0(n32930), .A1(n17694), .B0(n17072), .C0(n17071), .Y(
        n17073) );
  AOI211XL U21169 ( .A0(n17166), .A1(n17075), .B0(n17074), .C0(n17073), .Y(
        n17097) );
  AOI22XL U21170 ( .A0(n16744), .A1(weight_1[89]), .B0(weight_1[131]), .B1(
        n17801), .Y(n17079) );
  AOI22XL U21171 ( .A0(weight_1[167]), .A1(n17863), .B0(weight_1[77]), .B1(
        n17865), .Y(n17078) );
  AOI22XL U21172 ( .A0(weight_1[305]), .A1(n17798), .B0(weight_1[71]), .B1(
        n17883), .Y(n17077) );
  AOI22XL U21173 ( .A0(weight_1[221]), .A1(n17804), .B0(weight_1[113]), .B1(
        n17887), .Y(n17076) );
  NAND4XL U21174 ( .A(n17079), .B(n17078), .C(n17077), .D(n17076), .Y(n17095)
         );
  AOI22XL U21175 ( .A0(weight_1[311]), .A1(n17787), .B0(weight_1[143]), .B1(
        n17894), .Y(n17083) );
  AOI22XL U21176 ( .A0(weight_1[197]), .A1(n17866), .B0(weight_1[179]), .B1(
        n17899), .Y(n17082) );
  AOI22XL U21177 ( .A0(weight_1[53]), .A1(n17803), .B0(weight_1[29]), .B1(
        n17893), .Y(n17081) );
  AOI22XL U21178 ( .A0(weight_1[263]), .A1(n17886), .B0(weight_1[215]), .B1(
        n17898), .Y(n17080) );
  NAND4XL U21179 ( .A(n17083), .B(n17082), .C(n17081), .D(n17080), .Y(n17094)
         );
  AOI22XL U21180 ( .A0(n21766), .A1(weight_1[323]), .B0(weight_1[251]), .B1(
        n17797), .Y(n17087) );
  AOI22XL U21181 ( .A0(weight_1[395]), .A1(n17800), .B0(weight_1[161]), .B1(
        n17868), .Y(n17086) );
  AOI22XL U21182 ( .A0(weight_1[137]), .A1(n17895), .B0(weight_1[83]), .B1(
        n17799), .Y(n17085) );
  AOI22XL U21183 ( .A0(weight_1[149]), .A1(n17875), .B0(weight_1[41]), .B1(
        n17867), .Y(n17084) );
  NAND4XL U21184 ( .A(n17087), .B(n17086), .C(n17085), .D(n17084), .Y(n17093)
         );
  AOI22XL U21185 ( .A0(weight_1[281]), .A1(n17877), .B0(weight_1[227]), .B1(
        n17878), .Y(n17091) );
  AOI22XL U21186 ( .A0(weight_1[257]), .A1(n17896), .B0(weight_1[191]), .B1(
        n17790), .Y(n17090) );
  AOI22XL U21187 ( .A0(n21748), .A1(weight_1[317]), .B0(weight_1[35]), .B1(
        n17873), .Y(n17089) );
  AOI22XL U21188 ( .A0(n26082), .A1(weight_1[329]), .B0(weight_1[65]), .B1(
        n17791), .Y(n17088) );
  NAND4XL U21189 ( .A(n17091), .B(n17090), .C(n17089), .D(n17088), .Y(n17092)
         );
  NOR4XL U21190 ( .A(n17095), .B(n17094), .C(n17093), .D(n17092), .Y(n17096)
         );
  AOI32XL U21191 ( .A0(n17098), .A1(n17097), .A2(n17096), .B0(cursor[6]), .B1(
        n17097), .Y(n33404) );
  NAND2XL U21192 ( .A(n33404), .B(n20648), .Y(DP_OP_5166J1_122_9881_n70) );
  AOI22XL U21193 ( .A0(weight_1[463]), .A1(n17852), .B0(weight_1[457]), .B1(
        n17753), .Y(n17155) );
  AOI22XL U21194 ( .A0(weight_1[475]), .A1(n17842), .B0(weight_1[469]), .B1(
        n17691), .Y(n17154) );
  INVXL U21195 ( .A(weight_1[451]), .Y(n31328) );
  INVXL U21196 ( .A(weight_1[445]), .Y(n32727) );
  OAI22XL U21197 ( .A0(n31328), .A1(n17746), .B0(n32727), .B1(n17690), .Y(
        n17152) );
  AOI22XL U21198 ( .A0(weight_1[265]), .A1(n17788), .B0(weight_1[253]), .B1(
        n17896), .Y(n17102) );
  AOI22XL U21199 ( .A0(weight_1[187]), .A1(n17790), .B0(weight_1[25]), .B1(
        n17893), .Y(n17101) );
  AOI22XL U21200 ( .A0(n21999), .A1(weight_1[91]), .B0(weight_1[67]), .B1(
        n17883), .Y(n17100) );
  AOI22XL U21201 ( .A0(n21764), .A1(weight_1[19]), .B0(weight_1[169]), .B1(
        n17888), .Y(n17099) );
  NAND4XL U21202 ( .A(n17102), .B(n17101), .C(n17100), .D(n17099), .Y(n17118)
         );
  AOI22XL U21203 ( .A0(n26082), .A1(weight_1[325]), .B0(weight_1[73]), .B1(
        n17865), .Y(n17106) );
  AOI22XL U21204 ( .A0(n26059), .A1(weight_1[331]), .B0(weight_1[31]), .B1(
        n17873), .Y(n17105) );
  AOI22XL U21205 ( .A0(weight_1[211]), .A1(n17898), .B0(weight_1[79]), .B1(
        n17799), .Y(n17104) );
  AOI22XL U21206 ( .A0(weight_1[259]), .A1(n17886), .B0(weight_1[109]), .B1(
        n17887), .Y(n17103) );
  NAND4XL U21207 ( .A(n17106), .B(n17105), .C(n17104), .D(n17103), .Y(n17117)
         );
  AOI22XL U21208 ( .A0(weight_1[385]), .A1(n17821), .B0(weight_1[199]), .B1(
        n17813), .Y(n17110) );
  AOI22XL U21209 ( .A0(weight_1[379]), .A1(n17810), .B0(weight_1[337]), .B1(
        n17814), .Y(n17109) );
  AOI22XL U21210 ( .A0(weight_1[295]), .A1(n17826), .B0(weight_1[241]), .B1(
        n17815), .Y(n17108) );
  AOI22XL U21211 ( .A0(weight_1[349]), .A1(n17812), .B0(weight_1[235]), .B1(
        n17824), .Y(n17107) );
  NAND4XL U21212 ( .A(n17110), .B(n17109), .C(n17108), .D(n17107), .Y(n17116)
         );
  AOI22XL U21213 ( .A0(weight_1[343]), .A1(n17823), .B0(weight_1[133]), .B1(
        n17895), .Y(n17114) );
  AOI22XL U21214 ( .A0(weight_1[361]), .A1(n17827), .B0(weight_1[229]), .B1(
        n17811), .Y(n17113) );
  AOI22XL U21215 ( .A0(weight_1[373]), .A1(n17809), .B0(weight_1[367]), .B1(
        n17825), .Y(n17112) );
  AOI22XL U21216 ( .A0(weight_1[355]), .A1(n17816), .B0(weight_1[151]), .B1(
        n17822), .Y(n17111) );
  NAND4XL U21217 ( .A(n17114), .B(n17113), .C(n17112), .D(n17111), .Y(n17115)
         );
  AOI22XL U21218 ( .A0(weight_1[121]), .A1(n17792), .B0(weight_1[115]), .B1(
        n17876), .Y(n17122) );
  AOI22XL U21219 ( .A0(n21766), .A1(weight_1[319]), .B0(weight_1[247]), .B1(
        n17797), .Y(n17121) );
  AOI22XL U21220 ( .A0(weight_1[277]), .A1(n17877), .B0(weight_1[157]), .B1(
        n17868), .Y(n17120) );
  AOI22XL U21221 ( .A0(weight_1[205]), .A1(n17884), .B0(weight_1[175]), .B1(
        n17899), .Y(n17119) );
  NAND4XL U21222 ( .A(n17122), .B(n17121), .C(n17120), .D(n17119), .Y(n17138)
         );
  AOI22XL U21223 ( .A0(n21748), .A1(weight_1[313]), .B0(weight_1[49]), .B1(
        n17803), .Y(n17126) );
  AOI22XL U21224 ( .A0(weight_1[283]), .A1(n17802), .B0(weight_1[193]), .B1(
        n17866), .Y(n17125) );
  AOI22XL U21225 ( .A0(weight_1[163]), .A1(n17863), .B0(weight_1[97]), .B1(
        n17897), .Y(n17124) );
  AOI22XL U21226 ( .A0(weight_1[217]), .A1(n17804), .B0(weight_1[103]), .B1(
        n17885), .Y(n17123) );
  NAND4XL U21227 ( .A(n17126), .B(n17125), .C(n17124), .D(n17123), .Y(n17137)
         );
  AOI22XL U21228 ( .A0(n16744), .A1(weight_1[85]), .B0(weight_1[223]), .B1(
        n17878), .Y(n17130) );
  AOI22XL U21229 ( .A0(weight_1[145]), .A1(n17875), .B0(weight_1[55]), .B1(
        n17789), .Y(n17129) );
  AOI22XL U21230 ( .A0(weight_1[301]), .A1(n17798), .B0(weight_1[139]), .B1(
        n17894), .Y(n17128) );
  AOI22XL U21231 ( .A0(weight_1[127]), .A1(n17801), .B0(weight_1[61]), .B1(
        n17791), .Y(n17127) );
  NAND4XL U21232 ( .A(n17130), .B(n17129), .C(n17128), .D(n17127), .Y(n17136)
         );
  AOI22XL U21233 ( .A0(weight_1[391]), .A1(n17800), .B0(weight_1[307]), .B1(
        n17787), .Y(n17134) );
  AOI22XL U21234 ( .A0(weight_1[271]), .A1(n17864), .B0(weight_1[181]), .B1(
        n16724), .Y(n17133) );
  AOI22XL U21235 ( .A0(n21762), .A1(weight_1[13]), .B0(weight_1[289]), .B1(
        n17900), .Y(n17132) );
  AOI22XL U21236 ( .A0(weight_1[43]), .A1(n17874), .B0(weight_1[37]), .B1(
        n17867), .Y(n17131) );
  NAND4XL U21237 ( .A(n17134), .B(n17133), .C(n17132), .D(n17131), .Y(n17135)
         );
  AOI22XL U21238 ( .A0(n22021), .A1(weight_1[409]), .B0(n21887), .B1(
        weight_1[415]), .Y(n17142) );
  AOI22XL U21239 ( .A0(n16734), .A1(weight_1[403]), .B0(n21954), .B1(
        weight_1[397]), .Y(n17141) );
  AOI22XL U21240 ( .A0(n19475), .A1(weight_1[421]), .B0(n19097), .B1(
        weight_1[433]), .Y(n17140) );
  AOI22XL U21241 ( .A0(n19098), .A1(weight_1[439]), .B0(n19099), .B1(
        weight_1[427]), .Y(n17139) );
  NAND4XL U21242 ( .A(n17142), .B(n17141), .C(n17140), .D(n17139), .Y(n17147)
         );
  INVXL U21243 ( .A(weight_1[481]), .Y(n32415) );
  INVXL U21244 ( .A(weight_1[193]), .Y(n32496) );
  OAI22XL U21245 ( .A0(n17144), .A1(n32415), .B0(n32496), .B1(n17143), .Y(
        n17146) );
  INVXL U21246 ( .A(weight_1[391]), .Y(n32427) );
  INVXL U21247 ( .A(weight_1[1]), .Y(n32351) );
  OAI22XL U21248 ( .A0(n32427), .A1(n17391), .B0(n32351), .B1(n17188), .Y(
        n17145) );
  AOI211XL U21249 ( .A0(n16755), .A1(n17147), .B0(n17146), .C0(n17145), .Y(
        n17148) );
  AOI32XL U21250 ( .A0(n17150), .A1(n19182), .A2(n17149), .B0(cursor[6]), .B1(
        n17148), .Y(n17151) );
  AOI211XL U21251 ( .A0(weight_1[7]), .A1(n17444), .B0(n17152), .C0(n17151), 
        .Y(n17153) );
  NAND3X1 U21252 ( .A(n17155), .B(n17154), .C(n17153), .Y(n20619) );
  NAND2XL U21253 ( .A(n33554), .B(n20619), .Y(DP_OP_5166J1_122_9881_n56) );
  NAND2XL U21254 ( .A(n33404), .B(n20645), .Y(DP_OP_5166J1_122_9881_n76) );
  NAND2XL U21255 ( .A(n33554), .B(n17161), .Y(DP_OP_5166J1_122_9881_n54) );
  NAND2XL U21256 ( .A(n33554), .B(n20613), .Y(DP_OP_5166J1_122_9881_n55) );
  NAND2XL U21257 ( .A(n33404), .B(n17918), .Y(DP_OP_5166J1_122_9881_n58) );
  NAND2XL U21258 ( .A(n33554), .B(n17162), .Y(DP_OP_5166J1_122_9881_n53) );
  INVXL U21259 ( .A(affine_1[25]), .Y(DP_OP_5166J1_122_9881_n33) );
  AND2XL U21260 ( .A(n20619), .B(n20646), .Y(n17156) );
  AND2XL U21261 ( .A(n20619), .B(n17918), .Y(n17159) );
  AND2XL U21262 ( .A(n17161), .B(n20648), .Y(n17158) );
  ADDHXL U21263 ( .A(affine_1[23]), .B(n17156), .CO(n17157), .S(
        DP_OP_5166J1_122_9881_n45) );
  AND2XL U21264 ( .A(n20645), .B(n17161), .Y(DP_OP_5166J1_122_9881_n78) );
  AND2XL U21265 ( .A(n17162), .B(n20648), .Y(DP_OP_5166J1_122_9881_n71) );
  AND2XL U21266 ( .A(n17162), .B(n17918), .Y(n17164) );
  NAND2XL U21267 ( .A(n33404), .B(n20646), .Y(n17163) );
  AOI22XL U21268 ( .A0(weight_1[418]), .A1(n17854), .B0(weight_1[196]), .B1(
        n17813), .Y(n17225) );
  AOI22XL U21269 ( .A0(weight_1[472]), .A1(n17842), .B0(weight_1[466]), .B1(
        n17691), .Y(n17224) );
  INVXL U21270 ( .A(weight_1[442]), .Y(n32384) );
  OAI22XL U21271 ( .A0(n32385), .A1(n17746), .B0(n32384), .B1(n17690), .Y(
        n17179) );
  AOI22XL U21272 ( .A0(weight_1[436]), .A1(n17752), .B0(weight_1[430]), .B1(
        n17755), .Y(n17168) );
  NAND2XL U21273 ( .A(n21990), .B(n17166), .Y(n17748) );
  AOI22XL U21274 ( .A0(weight_1[412]), .A1(n17840), .B0(weight_1[406]), .B1(
        n17851), .Y(n17167) );
  OAI211XL U21275 ( .A0(n32910), .A1(n17248), .B0(n17168), .C0(n17167), .Y(
        n17178) );
  NAND2XL U21276 ( .A(n19097), .B(n17169), .Y(n17749) );
  OAI22XL U21277 ( .A0(n32759), .A1(n17749), .B0(n32386), .B1(n17837), .Y(
        n17177) );
  NOR2X2 U21278 ( .A(n26575), .B(n17170), .Y(n21752) );
  INVXL U21279 ( .A(n21752), .Y(n17171) );
  AOI21XL U21280 ( .A0(n17841), .A1(n18043), .B0(n17843), .Y(n17451) );
  INVXL U21281 ( .A(weight_1[484]), .Y(n32387) );
  AOI22XL U21282 ( .A0(weight_1[400]), .A1(n17853), .B0(weight_1[394]), .B1(
        n17754), .Y(n17175) );
  AOI22XL U21283 ( .A0(weight_1[460]), .A1(n17852), .B0(weight_1[424]), .B1(
        n17847), .Y(n17174) );
  OAI211XL U21284 ( .A0(n17451), .A1(n32387), .B0(n17175), .C0(n17174), .Y(
        n17176) );
  NOR4XL U21285 ( .A(n17179), .B(n17178), .C(n17177), .D(n17176), .Y(n17223)
         );
  AOI22XL U21286 ( .A0(weight_1[202]), .A1(n17884), .B0(weight_1[142]), .B1(
        n17875), .Y(n17183) );
  AOI22XL U21287 ( .A0(n21999), .A1(weight_1[88]), .B0(weight_1[256]), .B1(
        n17886), .Y(n17182) );
  AOI22XL U21288 ( .A0(weight_1[166]), .A1(n17888), .B0(weight_1[52]), .B1(
        n17789), .Y(n17181) );
  AOI22XL U21289 ( .A0(n21766), .A1(weight_1[316]), .B0(weight_1[190]), .B1(
        n17866), .Y(n17180) );
  NAND4XL U21290 ( .A(n17183), .B(n17182), .C(n17181), .D(n17180), .Y(n17221)
         );
  AOI22XL U21291 ( .A0(n26082), .A1(weight_1[322]), .B0(weight_1[214]), .B1(
        n17804), .Y(n17187) );
  AOI22XL U21292 ( .A0(weight_1[136]), .A1(n17894), .B0(weight_1[40]), .B1(
        n17874), .Y(n17186) );
  AOI22XL U21293 ( .A0(weight_1[274]), .A1(n17877), .B0(weight_1[22]), .B1(
        n17893), .Y(n17185) );
  AOI22XL U21294 ( .A0(n21764), .A1(weight_1[16]), .B0(weight_1[178]), .B1(
        n16724), .Y(n17184) );
  NAND4XL U21295 ( .A(n17187), .B(n17186), .C(n17185), .D(n17184), .Y(n17220)
         );
  AOI22XL U21296 ( .A0(weight_1[298]), .A1(n17798), .B0(weight_1[112]), .B1(
        n17876), .Y(n17218) );
  AOI22XL U21297 ( .A0(n16744), .A1(weight_1[82]), .B0(weight_1[280]), .B1(
        n17802), .Y(n17217) );
  INVXL U21298 ( .A(weight_1[10]), .Y(n32966) );
  INVXL U21299 ( .A(weight_1[382]), .Y(n32456) );
  OAI22XL U21300 ( .A0(n21556), .A1(n32966), .B0(n32456), .B1(n17188), .Y(
        n17194) );
  AOI22XL U21301 ( .A0(weight_1[262]), .A1(n17788), .B0(weight_1[100]), .B1(
        n17885), .Y(n17192) );
  AOI22XL U21302 ( .A0(weight_1[220]), .A1(n17878), .B0(weight_1[94]), .B1(
        n17897), .Y(n17191) );
  AOI22XL U21303 ( .A0(weight_1[244]), .A1(n17797), .B0(weight_1[106]), .B1(
        n17887), .Y(n17190) );
  AOI22XL U21304 ( .A0(weight_1[118]), .A1(n17792), .B0(weight_1[46]), .B1(
        n17803), .Y(n17189) );
  NAND4XL U21305 ( .A(n17192), .B(n17191), .C(n17190), .D(n17189), .Y(n17193)
         );
  AOI211XL U21306 ( .A0(weight_1[304]), .A1(n17787), .B0(n17194), .C0(n17193), 
        .Y(n17216) );
  AOI22XL U21307 ( .A0(weight_1[58]), .A1(n17791), .B0(weight_1[34]), .B1(
        n17867), .Y(n17198) );
  AOI22XL U21308 ( .A0(n21748), .A1(weight_1[310]), .B0(weight_1[124]), .B1(
        n17801), .Y(n17197) );
  AOI22XL U21309 ( .A0(n26059), .A1(weight_1[328]), .B0(weight_1[286]), .B1(
        n17900), .Y(n17196) );
  AOI22XL U21310 ( .A0(weight_1[130]), .A1(n17895), .B0(weight_1[70]), .B1(
        n17865), .Y(n17195) );
  NAND4XL U21311 ( .A(n17198), .B(n17197), .C(n17196), .D(n17195), .Y(n17214)
         );
  AOI22XL U21312 ( .A0(weight_1[388]), .A1(n17800), .B0(weight_1[64]), .B1(
        n17883), .Y(n17202) );
  AOI22XL U21313 ( .A0(weight_1[160]), .A1(n17863), .B0(weight_1[76]), .B1(
        n17799), .Y(n17201) );
  AOI22XL U21314 ( .A0(weight_1[268]), .A1(n17864), .B0(weight_1[250]), .B1(
        n17896), .Y(n17200) );
  AOI22XL U21315 ( .A0(weight_1[208]), .A1(n17898), .B0(weight_1[172]), .B1(
        n17899), .Y(n17199) );
  NAND4XL U21316 ( .A(n17202), .B(n17201), .C(n17200), .D(n17199), .Y(n17213)
         );
  AOI22XL U21317 ( .A0(weight_1[370]), .A1(n17809), .B0(weight_1[340]), .B1(
        n17823), .Y(n17206) );
  AOI22XL U21318 ( .A0(weight_1[376]), .A1(n17810), .B0(weight_1[148]), .B1(
        n17822), .Y(n17205) );
  AOI22XL U21319 ( .A0(weight_1[232]), .A1(n17824), .B0(weight_1[226]), .B1(
        n17811), .Y(n17204) );
  AOI22XL U21320 ( .A0(weight_1[358]), .A1(n17827), .B0(weight_1[352]), .B1(
        n17816), .Y(n17203) );
  NAND4XL U21321 ( .A(n17206), .B(n17205), .C(n17204), .D(n17203), .Y(n17212)
         );
  AOI22XL U21322 ( .A0(weight_1[184]), .A1(n17790), .B0(weight_1[154]), .B1(
        n17868), .Y(n17210) );
  AOI22XL U21323 ( .A0(weight_1[364]), .A1(n17825), .B0(weight_1[28]), .B1(
        n17873), .Y(n17209) );
  AOI22XL U21324 ( .A0(weight_1[346]), .A1(n17812), .B0(weight_1[292]), .B1(
        n17826), .Y(n17208) );
  AOI22XL U21325 ( .A0(weight_1[334]), .A1(n17814), .B0(weight_1[238]), .B1(
        n17815), .Y(n17207) );
  NAND4XL U21326 ( .A(n17210), .B(n17209), .C(n17208), .D(n17207), .Y(n17211)
         );
  NOR4XL U21327 ( .A(n17214), .B(n17213), .C(n17212), .D(n17211), .Y(n17215)
         );
  NAND4XL U21328 ( .A(n17218), .B(n17217), .C(n17216), .D(n17215), .Y(n17219)
         );
  OAI31XL U21329 ( .A0(n17221), .A1(n17220), .A2(n17219), .B0(n19182), .Y(
        n17222) );
  NAND4XL U21330 ( .A(n17225), .B(n17224), .C(n17223), .D(n17222), .Y(n17507)
         );
  NAND2XL U21331 ( .A(n20645), .B(n17507), .Y(n17505) );
  NAND2BXL U21332 ( .AN(affine_1[14]), .B(n17505), .Y(
        DP_OP_5167J1_123_9881_n39) );
  AOI22XL U21333 ( .A0(weight_1[201]), .A1(n17884), .B0(weight_1[171]), .B1(
        n17899), .Y(n17229) );
  AOI22XL U21334 ( .A0(n21748), .A1(weight_1[309]), .B0(weight_1[255]), .B1(
        n17886), .Y(n17228) );
  AOI22XL U21335 ( .A0(weight_1[273]), .A1(n17877), .B0(weight_1[117]), .B1(
        n17792), .Y(n17227) );
  AOI22XL U21336 ( .A0(weight_1[177]), .A1(n16724), .B0(weight_1[123]), .B1(
        n17801), .Y(n17226) );
  NAND4XL U21337 ( .A(n17229), .B(n17228), .C(n17227), .D(n17226), .Y(n17245)
         );
  AOI22XL U21338 ( .A0(n21766), .A1(weight_1[315]), .B0(weight_1[159]), .B1(
        n17863), .Y(n17233) );
  AOI22XL U21339 ( .A0(weight_1[267]), .A1(n17864), .B0(weight_1[243]), .B1(
        n17797), .Y(n17232) );
  AOI22XL U21340 ( .A0(weight_1[111]), .A1(n17876), .B0(weight_1[21]), .B1(
        n17893), .Y(n17231) );
  AOI22XL U21341 ( .A0(weight_1[249]), .A1(n17896), .B0(weight_1[207]), .B1(
        n17898), .Y(n17230) );
  NAND4XL U21342 ( .A(n17233), .B(n17232), .C(n17231), .D(n17230), .Y(n17244)
         );
  AOI22XL U21343 ( .A0(weight_1[333]), .A1(n17814), .B0(weight_1[225]), .B1(
        n17811), .Y(n17237) );
  AOI22XL U21344 ( .A0(weight_1[381]), .A1(n17821), .B0(weight_1[231]), .B1(
        n17824), .Y(n17236) );
  AOI22XL U21345 ( .A0(weight_1[357]), .A1(n17827), .B0(weight_1[345]), .B1(
        n17812), .Y(n17235) );
  AOI22XL U21346 ( .A0(weight_1[351]), .A1(n17816), .B0(weight_1[291]), .B1(
        n17826), .Y(n17234) );
  NAND4XL U21347 ( .A(n17237), .B(n17236), .C(n17235), .D(n17234), .Y(n17243)
         );
  AOI22XL U21348 ( .A0(weight_1[369]), .A1(n17809), .B0(weight_1[57]), .B1(
        n17791), .Y(n17241) );
  AOI22XL U21349 ( .A0(weight_1[363]), .A1(n17825), .B0(weight_1[195]), .B1(
        n17813), .Y(n17240) );
  AOI22XL U21350 ( .A0(weight_1[339]), .A1(n17823), .B0(weight_1[237]), .B1(
        n17815), .Y(n17239) );
  AOI22XL U21351 ( .A0(weight_1[375]), .A1(n17810), .B0(weight_1[147]), .B1(
        n17822), .Y(n17238) );
  NAND4XL U21352 ( .A(n17241), .B(n17240), .C(n17239), .D(n17238), .Y(n17242)
         );
  NOR4XL U21353 ( .A(n17245), .B(n17244), .C(n17243), .D(n17242), .Y(n17280)
         );
  INVXL U21354 ( .A(weight_1[3]), .Y(n32388) );
  AOI22XL U21355 ( .A0(weight_1[459]), .A1(n17852), .B0(weight_1[417]), .B1(
        n17854), .Y(n17247) );
  AOI22XL U21356 ( .A0(weight_1[465]), .A1(n17691), .B0(weight_1[441]), .B1(
        n17848), .Y(n17246) );
  OAI211XL U21357 ( .A0(n32388), .A1(n17248), .B0(n17247), .C0(n17246), .Y(
        n17257) );
  AOI22XL U21358 ( .A0(weight_1[435]), .A1(n17752), .B0(weight_1[393]), .B1(
        n17754), .Y(n17252) );
  AOI22XL U21359 ( .A0(weight_1[429]), .A1(n17755), .B0(weight_1[411]), .B1(
        n17840), .Y(n17251) );
  AOI22XL U21360 ( .A0(weight_1[477]), .A1(n17850), .B0(weight_1[423]), .B1(
        n17847), .Y(n17250) );
  AOI22XL U21361 ( .A0(weight_1[447]), .A1(n17849), .B0(weight_1[405]), .B1(
        n17851), .Y(n17249) );
  NAND4XL U21362 ( .A(n17252), .B(n17251), .C(n17250), .D(n17249), .Y(n17256)
         );
  OAI2BB2XL U21363 ( .B0(n32483), .B1(n17837), .A0N(weight_1[399]), .A1N(
        n17853), .Y(n17255) );
  INVXL U21364 ( .A(weight_1[483]), .Y(n32463) );
  AOI22XL U21365 ( .A0(n21763), .A1(weight_1[471]), .B0(weight_1[195]), .B1(
        n17813), .Y(n17253) );
  OAI22XL U21366 ( .A0(n17451), .A1(n32463), .B0(n17253), .B1(n19182), .Y(
        n17254) );
  NOR4XL U21367 ( .A(n17257), .B(n17256), .C(n17255), .D(n17254), .Y(n17279)
         );
  AOI22XL U21368 ( .A0(n26082), .A1(weight_1[321]), .B0(weight_1[39]), .B1(
        n17874), .Y(n17261) );
  AOI22XL U21369 ( .A0(n26059), .A1(weight_1[327]), .B0(n16744), .B1(
        weight_1[81]), .Y(n17260) );
  AOI22XL U21370 ( .A0(weight_1[51]), .A1(n17789), .B0(weight_1[33]), .B1(
        n17867), .Y(n17259) );
  AOI22XL U21371 ( .A0(weight_1[219]), .A1(n17878), .B0(weight_1[141]), .B1(
        n17875), .Y(n17258) );
  NAND4XL U21372 ( .A(n17261), .B(n17260), .C(n17259), .D(n17258), .Y(n17277)
         );
  AOI22XL U21373 ( .A0(n21764), .A1(weight_1[15]), .B0(weight_1[99]), .B1(
        n17885), .Y(n17265) );
  AOI22XL U21374 ( .A0(weight_1[387]), .A1(n17800), .B0(weight_1[303]), .B1(
        n17787), .Y(n17264) );
  AOI22XL U21375 ( .A0(weight_1[285]), .A1(n17900), .B0(weight_1[45]), .B1(
        n17803), .Y(n17263) );
  AOI22XL U21376 ( .A0(n21762), .A1(weight_1[9]), .B0(weight_1[213]), .B1(
        n17804), .Y(n17262) );
  NAND4XL U21377 ( .A(n17265), .B(n17264), .C(n17263), .D(n17262), .Y(n17276)
         );
  AOI22XL U21378 ( .A0(weight_1[183]), .A1(n17790), .B0(weight_1[75]), .B1(
        n17799), .Y(n17269) );
  AOI22XL U21379 ( .A0(n21999), .A1(weight_1[87]), .B0(weight_1[261]), .B1(
        n17788), .Y(n17268) );
  AOI22XL U21380 ( .A0(weight_1[63]), .A1(n17883), .B0(weight_1[27]), .B1(
        n17873), .Y(n17267) );
  AOI22XL U21381 ( .A0(weight_1[135]), .A1(n17894), .B0(weight_1[93]), .B1(
        n17897), .Y(n17266) );
  NAND4XL U21382 ( .A(n17269), .B(n17268), .C(n17267), .D(n17266), .Y(n17275)
         );
  AOI22XL U21383 ( .A0(weight_1[153]), .A1(n17868), .B0(weight_1[105]), .B1(
        n17887), .Y(n17273) );
  AOI22XL U21384 ( .A0(weight_1[189]), .A1(n17866), .B0(weight_1[129]), .B1(
        n17895), .Y(n17272) );
  AOI22XL U21385 ( .A0(weight_1[297]), .A1(n17798), .B0(weight_1[165]), .B1(
        n17888), .Y(n17271) );
  AOI22XL U21386 ( .A0(weight_1[279]), .A1(n17802), .B0(weight_1[69]), .B1(
        n17865), .Y(n17270) );
  NAND4XL U21387 ( .A(n17273), .B(n17272), .C(n17271), .D(n17270), .Y(n17274)
         );
  NOR4XL U21388 ( .A(n17277), .B(n17276), .C(n17275), .D(n17274), .Y(n17278)
         );
  AOI32XL U21389 ( .A0(n17280), .A1(n17279), .A2(n17278), .B0(cursor[6]), .B1(
        n17279), .Y(n17506) );
  AND2XL U21390 ( .A(n17506), .B(n17918), .Y(DP_OP_5167J1_123_9881_n60) );
  AOI22XL U21391 ( .A0(weight_1[464]), .A1(n17691), .B0(weight_1[398]), .B1(
        n17853), .Y(n17334) );
  AOI22XL U21392 ( .A0(weight_1[194]), .A1(n17813), .B0(weight_1[2]), .B1(
        n17444), .Y(n17333) );
  INVXL U21393 ( .A(weight_1[452]), .Y(n32379) );
  INVXL U21394 ( .A(weight_1[404]), .Y(n32733) );
  OAI22XL U21395 ( .A0(n32379), .A1(n17837), .B0(n32733), .B1(n17748), .Y(
        n17288) );
  INVXL U21396 ( .A(weight_1[470]), .Y(n32355) );
  AOI22XL U21397 ( .A0(weight_1[410]), .A1(n17840), .B0(weight_1[392]), .B1(
        n17754), .Y(n17282) );
  AOI22XL U21398 ( .A0(weight_1[476]), .A1(n17850), .B0(weight_1[416]), .B1(
        n17854), .Y(n17281) );
  OAI211XL U21399 ( .A0(n32355), .A1(n17694), .B0(n17282), .C0(n17281), .Y(
        n17287) );
  INVXL U21400 ( .A(weight_1[446]), .Y(n32380) );
  INVXL U21401 ( .A(weight_1[440]), .Y(n32375) );
  OAI22XL U21402 ( .A0(n32380), .A1(n17746), .B0(n32375), .B1(n17690), .Y(
        n17286) );
  INVXL U21403 ( .A(weight_1[482]), .Y(n32678) );
  AOI22XL U21404 ( .A0(weight_1[434]), .A1(n17752), .B0(weight_1[422]), .B1(
        n17847), .Y(n17284) );
  AOI22XL U21405 ( .A0(weight_1[458]), .A1(n17852), .B0(weight_1[428]), .B1(
        n17755), .Y(n17283) );
  OAI211XL U21406 ( .A0(n17451), .A1(n32678), .B0(n17284), .C0(n17283), .Y(
        n17285) );
  NOR4XL U21407 ( .A(n17288), .B(n17287), .C(n17286), .D(n17285), .Y(n17332)
         );
  AOI22XL U21408 ( .A0(weight_1[248]), .A1(n17896), .B0(weight_1[134]), .B1(
        n17894), .Y(n17292) );
  AOI22XL U21409 ( .A0(weight_1[164]), .A1(n17888), .B0(weight_1[32]), .B1(
        n17867), .Y(n17291) );
  AOI22XL U21410 ( .A0(n21762), .A1(weight_1[8]), .B0(weight_1[128]), .B1(
        n17895), .Y(n17290) );
  AOI22XL U21411 ( .A0(weight_1[170]), .A1(n17899), .B0(weight_1[116]), .B1(
        n17792), .Y(n17289) );
  NAND4XL U21412 ( .A(n17292), .B(n17291), .C(n17290), .D(n17289), .Y(n17330)
         );
  AOI22XL U21413 ( .A0(weight_1[302]), .A1(n17787), .B0(weight_1[212]), .B1(
        n17804), .Y(n17296) );
  AOI22XL U21414 ( .A0(n21999), .A1(weight_1[86]), .B0(weight_1[266]), .B1(
        n17864), .Y(n17295) );
  AOI22XL U21415 ( .A0(weight_1[74]), .A1(n17799), .B0(weight_1[56]), .B1(
        n17791), .Y(n17294) );
  AOI22XL U21416 ( .A0(n21766), .A1(weight_1[314]), .B0(weight_1[188]), .B1(
        n17866), .Y(n17293) );
  NAND4XL U21417 ( .A(n17296), .B(n17295), .C(n17294), .D(n17293), .Y(n17329)
         );
  AOI22XL U21418 ( .A0(n26059), .A1(weight_1[326]), .B0(weight_1[284]), .B1(
        n17900), .Y(n17327) );
  AOI22XL U21419 ( .A0(weight_1[104]), .A1(n17887), .B0(weight_1[38]), .B1(
        n17874), .Y(n17326) );
  AOI22XL U21420 ( .A0(weight_1[110]), .A1(n17876), .B0(weight_1[68]), .B1(
        n17865), .Y(n17297) );
  INVXL U21421 ( .A(n17297), .Y(n17303) );
  AOI22XL U21422 ( .A0(n26082), .A1(weight_1[320]), .B0(weight_1[98]), .B1(
        n17885), .Y(n17301) );
  AOI22XL U21423 ( .A0(weight_1[200]), .A1(n17884), .B0(weight_1[44]), .B1(
        n17803), .Y(n17300) );
  AOI22XL U21424 ( .A0(weight_1[242]), .A1(n17797), .B0(weight_1[92]), .B1(
        n17897), .Y(n17299) );
  AOI22XL U21425 ( .A0(weight_1[386]), .A1(n17800), .B0(weight_1[152]), .B1(
        n17868), .Y(n17298) );
  NAND4XL U21426 ( .A(n17301), .B(n17300), .C(n17299), .D(n17298), .Y(n17302)
         );
  AOI211XL U21427 ( .A0(weight_1[236]), .A1(n17815), .B0(n17303), .C0(n17302), 
        .Y(n17325) );
  AOI22XL U21428 ( .A0(n21748), .A1(weight_1[308]), .B0(weight_1[176]), .B1(
        n16724), .Y(n17307) );
  AOI22XL U21429 ( .A0(weight_1[140]), .A1(n17875), .B0(weight_1[26]), .B1(
        n17873), .Y(n17306) );
  AOI22XL U21430 ( .A0(n16744), .A1(weight_1[80]), .B0(weight_1[206]), .B1(
        n17898), .Y(n17305) );
  AOI22XL U21431 ( .A0(weight_1[218]), .A1(n17878), .B0(weight_1[158]), .B1(
        n17863), .Y(n17304) );
  NAND4XL U21432 ( .A(n17307), .B(n17306), .C(n17305), .D(n17304), .Y(n17323)
         );
  AOI22XL U21433 ( .A0(weight_1[254]), .A1(n17886), .B0(weight_1[182]), .B1(
        n17790), .Y(n17311) );
  AOI22XL U21434 ( .A0(weight_1[278]), .A1(n17802), .B0(weight_1[260]), .B1(
        n17788), .Y(n17310) );
  AOI22XL U21435 ( .A0(weight_1[272]), .A1(n17877), .B0(weight_1[62]), .B1(
        n17883), .Y(n17309) );
  AOI22XL U21436 ( .A0(weight_1[296]), .A1(n17798), .B0(weight_1[122]), .B1(
        n17801), .Y(n17308) );
  NAND4XL U21437 ( .A(n17311), .B(n17310), .C(n17309), .D(n17308), .Y(n17322)
         );
  AOI22XL U21438 ( .A0(weight_1[332]), .A1(n17814), .B0(weight_1[224]), .B1(
        n17811), .Y(n17315) );
  AOI22XL U21439 ( .A0(weight_1[230]), .A1(n17824), .B0(weight_1[146]), .B1(
        n17822), .Y(n17314) );
  AOI22XL U21440 ( .A0(weight_1[374]), .A1(n17810), .B0(weight_1[290]), .B1(
        n17826), .Y(n17313) );
  AOI22XL U21441 ( .A0(weight_1[350]), .A1(n17816), .B0(weight_1[338]), .B1(
        n17823), .Y(n17312) );
  NAND4XL U21442 ( .A(n17315), .B(n17314), .C(n17313), .D(n17312), .Y(n17321)
         );
  AOI22XL U21443 ( .A0(n21764), .A1(weight_1[14]), .B0(weight_1[50]), .B1(
        n17789), .Y(n17319) );
  AOI22XL U21444 ( .A0(weight_1[356]), .A1(n17827), .B0(weight_1[20]), .B1(
        n17893), .Y(n17318) );
  AOI22XL U21445 ( .A0(weight_1[362]), .A1(n17825), .B0(weight_1[344]), .B1(
        n17812), .Y(n17317) );
  AOI22XL U21446 ( .A0(weight_1[380]), .A1(n17821), .B0(weight_1[368]), .B1(
        n17809), .Y(n17316) );
  NAND4XL U21447 ( .A(n17319), .B(n17318), .C(n17317), .D(n17316), .Y(n17320)
         );
  NOR4XL U21448 ( .A(n17323), .B(n17322), .C(n17321), .D(n17320), .Y(n17324)
         );
  NAND4XL U21449 ( .A(n17327), .B(n17326), .C(n17325), .D(n17324), .Y(n17328)
         );
  OAI31XL U21450 ( .A0(n17330), .A1(n17329), .A2(n17328), .B0(n19182), .Y(
        n17331) );
  NAND4XL U21451 ( .A(n17334), .B(n17333), .C(n17332), .D(n17331), .Y(n20628)
         );
  AND2XL U21452 ( .A(n20628), .B(n17918), .Y(DP_OP_5167J1_123_9881_n61) );
  AND2XL U21453 ( .A(n17507), .B(n20646), .Y(DP_OP_5167J1_123_9881_n65) );
  AND2XL U21454 ( .A(n20628), .B(n20646), .Y(DP_OP_5167J1_123_9881_n67) );
  AND2XL U21455 ( .A(n20628), .B(n20648), .Y(DP_OP_5167J1_123_9881_n73) );
  AOI22XL U21456 ( .A0(weight_1[473]), .A1(n17842), .B0(weight_1[413]), .B1(
        n17840), .Y(n17388) );
  AOI22XL U21457 ( .A0(weight_1[467]), .A1(n17691), .B0(weight_1[5]), .B1(
        n17444), .Y(n17387) );
  AOI22XL U21458 ( .A0(weight_1[449]), .A1(n17849), .B0(weight_1[443]), .B1(
        n17848), .Y(n17338) );
  AOI22XL U21459 ( .A0(weight_1[461]), .A1(n17852), .B0(weight_1[395]), .B1(
        n17754), .Y(n17337) );
  AOI22XL U21460 ( .A0(weight_1[455]), .A1(n17753), .B0(weight_1[425]), .B1(
        n17847), .Y(n17336) );
  AOI22XL U21461 ( .A0(weight_1[437]), .A1(n17752), .B0(weight_1[407]), .B1(
        n17851), .Y(n17335) );
  NAND4XL U21462 ( .A(n17338), .B(n17337), .C(n17336), .D(n17335), .Y(n17342)
         );
  INVXL U21463 ( .A(weight_1[485]), .Y(n32929) );
  AOI22XL U21464 ( .A0(weight_1[479]), .A1(n17850), .B0(weight_1[419]), .B1(
        n17854), .Y(n17340) );
  AOI22XL U21465 ( .A0(weight_1[431]), .A1(n17755), .B0(weight_1[401]), .B1(
        n17853), .Y(n17339) );
  OAI211XL U21466 ( .A0(n17451), .A1(n32929), .B0(n17340), .C0(n17339), .Y(
        n17341) );
  AOI211XL U21467 ( .A0(weight_1[197]), .A1(n17454), .B0(n17342), .C0(n17341), 
        .Y(n17386) );
  AOI22XL U21468 ( .A0(weight_1[47]), .A1(n17803), .B0(weight_1[29]), .B1(
        n17873), .Y(n17346) );
  AOI22XL U21469 ( .A0(weight_1[305]), .A1(n17787), .B0(weight_1[35]), .B1(
        n17867), .Y(n17345) );
  AOI22XL U21470 ( .A0(weight_1[95]), .A1(n17897), .B0(weight_1[53]), .B1(
        n17789), .Y(n17344) );
  AOI22XL U21471 ( .A0(weight_1[281]), .A1(n17802), .B0(weight_1[155]), .B1(
        n17868), .Y(n17343) );
  NAND4XL U21472 ( .A(n17346), .B(n17345), .C(n17344), .D(n17343), .Y(n17362)
         );
  AOI22XL U21473 ( .A0(weight_1[125]), .A1(n17801), .B0(weight_1[65]), .B1(
        n17883), .Y(n17350) );
  AOI22XL U21474 ( .A0(n26082), .A1(weight_1[323]), .B0(weight_1[131]), .B1(
        n17895), .Y(n17349) );
  AOI22XL U21475 ( .A0(weight_1[113]), .A1(n17876), .B0(weight_1[23]), .B1(
        n17893), .Y(n17348) );
  AOI22XL U21476 ( .A0(weight_1[287]), .A1(n17900), .B0(weight_1[161]), .B1(
        n17863), .Y(n17347) );
  NAND4XL U21477 ( .A(n17350), .B(n17349), .C(n17348), .D(n17347), .Y(n17361)
         );
  AOI22XL U21478 ( .A0(weight_1[359]), .A1(n17827), .B0(weight_1[341]), .B1(
        n17823), .Y(n17354) );
  AOI22XL U21479 ( .A0(weight_1[293]), .A1(n17826), .B0(weight_1[233]), .B1(
        n17824), .Y(n17353) );
  AOI22XL U21480 ( .A0(weight_1[353]), .A1(n17816), .B0(weight_1[347]), .B1(
        n17812), .Y(n17352) );
  AOI22XL U21481 ( .A0(weight_1[377]), .A1(n17810), .B0(weight_1[197]), .B1(
        n17813), .Y(n17351) );
  NAND4XL U21482 ( .A(n17354), .B(n17353), .C(n17352), .D(n17351), .Y(n17360)
         );
  AOI22XL U21483 ( .A0(weight_1[239]), .A1(n17815), .B0(weight_1[71]), .B1(
        n17865), .Y(n17358) );
  AOI22XL U21484 ( .A0(weight_1[383]), .A1(n17821), .B0(weight_1[227]), .B1(
        n17811), .Y(n17357) );
  AOI22XL U21485 ( .A0(weight_1[365]), .A1(n17825), .B0(weight_1[335]), .B1(
        n17814), .Y(n17356) );
  AOI22XL U21486 ( .A0(weight_1[371]), .A1(n17809), .B0(weight_1[149]), .B1(
        n17822), .Y(n17355) );
  NAND4XL U21487 ( .A(n17358), .B(n17357), .C(n17356), .D(n17355), .Y(n17359)
         );
  NOR4XL U21488 ( .A(n17362), .B(n17361), .C(n17360), .D(n17359), .Y(n17384)
         );
  AOI22XL U21489 ( .A0(n21764), .A1(weight_1[17]), .B0(weight_1[173]), .B1(
        n17899), .Y(n17366) );
  AOI22XL U21490 ( .A0(weight_1[263]), .A1(n17788), .B0(weight_1[215]), .B1(
        n17804), .Y(n17365) );
  AOI22XL U21491 ( .A0(weight_1[209]), .A1(n17898), .B0(weight_1[203]), .B1(
        n17884), .Y(n17364) );
  AOI22XL U21492 ( .A0(n16744), .A1(weight_1[83]), .B0(weight_1[275]), .B1(
        n17877), .Y(n17363) );
  NAND4XL U21493 ( .A(n17366), .B(n17365), .C(n17364), .D(n17363), .Y(n17382)
         );
  AOI22XL U21494 ( .A0(weight_1[299]), .A1(n17798), .B0(weight_1[269]), .B1(
        n17864), .Y(n17370) );
  AOI22XL U21495 ( .A0(n21999), .A1(weight_1[89]), .B0(weight_1[101]), .B1(
        n17885), .Y(n17369) );
  AOI22XL U21496 ( .A0(weight_1[179]), .A1(n16724), .B0(weight_1[77]), .B1(
        n17799), .Y(n17368) );
  AOI22XL U21497 ( .A0(weight_1[257]), .A1(n17886), .B0(weight_1[119]), .B1(
        n17792), .Y(n17367) );
  NAND4XL U21498 ( .A(n17370), .B(n17369), .C(n17368), .D(n17367), .Y(n17381)
         );
  AOI22XL U21499 ( .A0(n26059), .A1(weight_1[329]), .B0(weight_1[107]), .B1(
        n17887), .Y(n17374) );
  AOI22XL U21500 ( .A0(weight_1[137]), .A1(n17894), .B0(weight_1[41]), .B1(
        n17874), .Y(n17373) );
  AOI22XL U21501 ( .A0(weight_1[245]), .A1(n17797), .B0(weight_1[143]), .B1(
        n17875), .Y(n17372) );
  AOI22XL U21502 ( .A0(n21766), .A1(weight_1[317]), .B0(weight_1[221]), .B1(
        n17878), .Y(n17371) );
  NAND4XL U21503 ( .A(n17374), .B(n17373), .C(n17372), .D(n17371), .Y(n17380)
         );
  AOI22XL U21504 ( .A0(weight_1[185]), .A1(n17790), .B0(weight_1[59]), .B1(
        n17791), .Y(n17378) );
  AOI22XL U21505 ( .A0(weight_1[389]), .A1(n17800), .B0(weight_1[251]), .B1(
        n17896), .Y(n17377) );
  AOI22XL U21506 ( .A0(n21762), .A1(weight_1[11]), .B0(weight_1[191]), .B1(
        n17866), .Y(n17376) );
  AOI22XL U21507 ( .A0(n21748), .A1(weight_1[311]), .B0(weight_1[167]), .B1(
        n17888), .Y(n17375) );
  NAND4XL U21508 ( .A(n17378), .B(n17377), .C(n17376), .D(n17375), .Y(n17379)
         );
  NOR4XL U21509 ( .A(n17382), .B(n17381), .C(n17380), .D(n17379), .Y(n17383)
         );
  OAI2BB1XL U21510 ( .A0N(n17384), .A1N(n17383), .B0(n19182), .Y(n17385) );
  NAND4XL U21511 ( .A(n17388), .B(n17387), .C(n17386), .D(n17385), .Y(n33553)
         );
  NAND2XL U21512 ( .A(n33553), .B(n20648), .Y(DP_OP_5167J1_123_9881_n70) );
  AOI22XL U21513 ( .A0(weight_1[468]), .A1(n17842), .B0(weight_1[402]), .B1(
        n17851), .Y(n17443) );
  AOI22XL U21514 ( .A0(weight_1[462]), .A1(n17691), .B0(weight_1[0]), .B1(
        n17444), .Y(n17442) );
  INVXL U21515 ( .A(weight_1[474]), .Y(n26914) );
  INVXL U21516 ( .A(weight_1[390]), .Y(n26900) );
  INVXL U21517 ( .A(n17754), .Y(n17838) );
  OAI22XL U21518 ( .A0(n26914), .A1(n17749), .B0(n26900), .B1(n17838), .Y(
        n17397) );
  AOI22XL U21519 ( .A0(weight_1[432]), .A1(n17752), .B0(weight_1[396]), .B1(
        n17853), .Y(n17390) );
  AOI22XL U21520 ( .A0(weight_1[426]), .A1(n17755), .B0(weight_1[420]), .B1(
        n17847), .Y(n17389) );
  OAI211XL U21521 ( .A0(n26868), .A1(n17391), .B0(n17390), .C0(n17389), .Y(
        n17396) );
  INVXL U21522 ( .A(weight_1[444]), .Y(n26854) );
  OAI22XL U21523 ( .A0(n26854), .A1(n17746), .B0(n26885), .B1(n17690), .Y(
        n17395) );
  INVXL U21524 ( .A(weight_1[480]), .Y(n26913) );
  AOI22XL U21525 ( .A0(weight_1[456]), .A1(n17852), .B0(weight_1[408]), .B1(
        n17840), .Y(n17393) );
  AOI22XL U21526 ( .A0(weight_1[450]), .A1(n17753), .B0(weight_1[414]), .B1(
        n17854), .Y(n17392) );
  OAI211XL U21527 ( .A0(n17451), .A1(n26913), .B0(n17393), .C0(n17392), .Y(
        n17394) );
  NOR4XL U21528 ( .A(n17397), .B(n17396), .C(n17395), .D(n17394), .Y(n17441)
         );
  AOI22XL U21529 ( .A0(weight_1[258]), .A1(n17788), .B0(weight_1[240]), .B1(
        n17797), .Y(n17401) );
  AOI22XL U21530 ( .A0(n21764), .A1(weight_1[12]), .B0(weight_1[42]), .B1(
        n17803), .Y(n17400) );
  AOI22XL U21531 ( .A0(weight_1[264]), .A1(n17864), .B0(weight_1[24]), .B1(
        n17873), .Y(n17399) );
  AOI22XL U21532 ( .A0(weight_1[150]), .A1(n17868), .B0(weight_1[96]), .B1(
        n17885), .Y(n17398) );
  NAND4XL U21533 ( .A(n17401), .B(n17400), .C(n17399), .D(n17398), .Y(n17439)
         );
  AOI22XL U21534 ( .A0(n21999), .A1(weight_1[84]), .B0(weight_1[174]), .B1(
        n16724), .Y(n17405) );
  AOI22XL U21535 ( .A0(n16744), .A1(weight_1[78]), .B0(n21748), .B1(
        weight_1[306]), .Y(n17404) );
  AOI22XL U21536 ( .A0(weight_1[276]), .A1(n17802), .B0(weight_1[156]), .B1(
        n17863), .Y(n17403) );
  AOI22XL U21537 ( .A0(weight_1[180]), .A1(n17790), .B0(weight_1[126]), .B1(
        n17895), .Y(n17402) );
  NAND4XL U21538 ( .A(n17405), .B(n17404), .C(n17403), .D(n17402), .Y(n17438)
         );
  AOI22XL U21539 ( .A0(weight_1[294]), .A1(n17798), .B0(weight_1[120]), .B1(
        n17801), .Y(n17436) );
  AOI22XL U21540 ( .A0(weight_1[270]), .A1(n17877), .B0(weight_1[186]), .B1(
        n17866), .Y(n17435) );
  AOI22XL U21541 ( .A0(weight_1[204]), .A1(n17898), .B0(weight_1[60]), .B1(
        n17883), .Y(n17406) );
  INVXL U21542 ( .A(n17406), .Y(n17412) );
  AOI22XL U21543 ( .A0(weight_1[132]), .A1(n17894), .B0(weight_1[18]), .B1(
        n17893), .Y(n17410) );
  AOI22XL U21544 ( .A0(weight_1[216]), .A1(n17878), .B0(weight_1[108]), .B1(
        n17876), .Y(n17409) );
  AOI22XL U21545 ( .A0(n26082), .A1(weight_1[318]), .B0(weight_1[90]), .B1(
        n17897), .Y(n17408) );
  AOI22XL U21546 ( .A0(n21762), .A1(weight_1[6]), .B0(weight_1[66]), .B1(
        n17865), .Y(n17407) );
  NAND4XL U21547 ( .A(n17410), .B(n17409), .C(n17408), .D(n17407), .Y(n17411)
         );
  AOI211XL U21548 ( .A0(weight_1[288]), .A1(n17826), .B0(n17412), .C0(n17411), 
        .Y(n17434) );
  AOI22XL U21549 ( .A0(weight_1[138]), .A1(n17875), .B0(weight_1[102]), .B1(
        n17887), .Y(n17416) );
  AOI22XL U21550 ( .A0(weight_1[252]), .A1(n17886), .B0(weight_1[72]), .B1(
        n17799), .Y(n17415) );
  AOI22XL U21551 ( .A0(n26059), .A1(weight_1[324]), .B0(weight_1[300]), .B1(
        n17787), .Y(n17414) );
  AOI22XL U21552 ( .A0(weight_1[282]), .A1(n17900), .B0(weight_1[30]), .B1(
        n17867), .Y(n17413) );
  NAND4XL U21553 ( .A(n17416), .B(n17415), .C(n17414), .D(n17413), .Y(n17432)
         );
  AOI22XL U21554 ( .A0(weight_1[246]), .A1(n17896), .B0(weight_1[54]), .B1(
        n17791), .Y(n17420) );
  AOI22XL U21555 ( .A0(weight_1[168]), .A1(n17899), .B0(weight_1[48]), .B1(
        n17789), .Y(n17419) );
  AOI22XL U21556 ( .A0(weight_1[384]), .A1(n17800), .B0(weight_1[210]), .B1(
        n17804), .Y(n17418) );
  AOI22XL U21557 ( .A0(n21766), .A1(weight_1[312]), .B0(weight_1[114]), .B1(
        n17792), .Y(n17417) );
  NAND4XL U21558 ( .A(n17420), .B(n17419), .C(n17418), .D(n17417), .Y(n17431)
         );
  AOI22XL U21559 ( .A0(weight_1[372]), .A1(n17810), .B0(weight_1[348]), .B1(
        n17816), .Y(n17424) );
  AOI22XL U21560 ( .A0(weight_1[360]), .A1(n17825), .B0(weight_1[222]), .B1(
        n17811), .Y(n17423) );
  AOI22XL U21561 ( .A0(weight_1[366]), .A1(n17809), .B0(weight_1[354]), .B1(
        n17827), .Y(n17422) );
  AOI22XL U21562 ( .A0(weight_1[342]), .A1(n17812), .B0(weight_1[336]), .B1(
        n17823), .Y(n17421) );
  NAND4XL U21563 ( .A(n17424), .B(n17423), .C(n17422), .D(n17421), .Y(n17430)
         );
  AOI22XL U21564 ( .A0(weight_1[198]), .A1(n17884), .B0(weight_1[162]), .B1(
        n17888), .Y(n17428) );
  AOI22XL U21565 ( .A0(weight_1[330]), .A1(n17814), .B0(weight_1[36]), .B1(
        n17874), .Y(n17427) );
  AOI22XL U21566 ( .A0(weight_1[228]), .A1(n17824), .B0(weight_1[144]), .B1(
        n17822), .Y(n17426) );
  AOI22XL U21567 ( .A0(weight_1[378]), .A1(n17821), .B0(weight_1[234]), .B1(
        n17815), .Y(n17425) );
  NAND4XL U21568 ( .A(n17428), .B(n17427), .C(n17426), .D(n17425), .Y(n17429)
         );
  NOR4XL U21569 ( .A(n17432), .B(n17431), .C(n17430), .D(n17429), .Y(n17433)
         );
  NAND2XL U21570 ( .A(n33554), .B(n20634), .Y(DP_OP_5167J1_123_9881_n57) );
  AOI22XL U21571 ( .A0(weight_1[475]), .A1(n17850), .B0(weight_1[469]), .B1(
        n17842), .Y(n17500) );
  AOI22XL U21572 ( .A0(weight_1[463]), .A1(n17691), .B0(weight_1[1]), .B1(
        n17444), .Y(n17499) );
  AOI22XL U21573 ( .A0(weight_1[433]), .A1(n17752), .B0(weight_1[421]), .B1(
        n17847), .Y(n17448) );
  AOI22XL U21574 ( .A0(weight_1[397]), .A1(n17853), .B0(weight_1[391]), .B1(
        n17754), .Y(n17447) );
  AOI22XL U21575 ( .A0(weight_1[457]), .A1(n17852), .B0(weight_1[415]), .B1(
        n17854), .Y(n17446) );
  AOI22XL U21576 ( .A0(weight_1[451]), .A1(n17753), .B0(weight_1[439]), .B1(
        n17848), .Y(n17445) );
  NAND4XL U21577 ( .A(n17448), .B(n17447), .C(n17446), .D(n17445), .Y(n17453)
         );
  AOI22XL U21578 ( .A0(weight_1[445]), .A1(n17849), .B0(weight_1[427]), .B1(
        n17755), .Y(n17450) );
  AOI22XL U21579 ( .A0(weight_1[409]), .A1(n17840), .B0(weight_1[403]), .B1(
        n17851), .Y(n17449) );
  OAI211XL U21580 ( .A0(n17451), .A1(n32415), .B0(n17450), .C0(n17449), .Y(
        n17452) );
  AOI211XL U21581 ( .A0(weight_1[193]), .A1(n17454), .B0(n17453), .C0(n17452), 
        .Y(n17498) );
  AOI22XL U21582 ( .A0(weight_1[253]), .A1(n17886), .B0(weight_1[217]), .B1(
        n17878), .Y(n17458) );
  AOI22XL U21583 ( .A0(weight_1[205]), .A1(n17898), .B0(weight_1[187]), .B1(
        n17866), .Y(n17457) );
  AOI22XL U21584 ( .A0(weight_1[169]), .A1(n17899), .B0(weight_1[133]), .B1(
        n17894), .Y(n17456) );
  AOI22XL U21585 ( .A0(weight_1[115]), .A1(n17792), .B0(weight_1[19]), .B1(
        n17893), .Y(n17455) );
  NAND4XL U21586 ( .A(n17458), .B(n17457), .C(n17456), .D(n17455), .Y(n17474)
         );
  AOI22XL U21587 ( .A0(n21999), .A1(weight_1[85]), .B0(weight_1[97]), .B1(
        n17885), .Y(n17462) );
  AOI22XL U21588 ( .A0(n26059), .A1(weight_1[325]), .B0(weight_1[283]), .B1(
        n17900), .Y(n17461) );
  AOI22XL U21589 ( .A0(weight_1[265]), .A1(n17864), .B0(weight_1[127]), .B1(
        n17895), .Y(n17460) );
  AOI22XL U21590 ( .A0(weight_1[211]), .A1(n17804), .B0(weight_1[175]), .B1(
        n16724), .Y(n17459) );
  NAND4XL U21591 ( .A(n17462), .B(n17461), .C(n17460), .D(n17459), .Y(n17473)
         );
  AOI22XL U21592 ( .A0(weight_1[361]), .A1(n17825), .B0(weight_1[337]), .B1(
        n17823), .Y(n17466) );
  AOI22XL U21593 ( .A0(weight_1[331]), .A1(n17814), .B0(weight_1[289]), .B1(
        n17826), .Y(n17465) );
  AOI22XL U21594 ( .A0(weight_1[343]), .A1(n17812), .B0(weight_1[193]), .B1(
        n17813), .Y(n17464) );
  AOI22XL U21595 ( .A0(weight_1[373]), .A1(n17810), .B0(weight_1[349]), .B1(
        n17816), .Y(n17463) );
  NAND4XL U21596 ( .A(n17466), .B(n17465), .C(n17464), .D(n17463), .Y(n17472)
         );
  AOI22XL U21597 ( .A0(weight_1[229]), .A1(n17824), .B0(weight_1[109]), .B1(
        n17876), .Y(n17470) );
  AOI22XL U21598 ( .A0(weight_1[367]), .A1(n17809), .B0(weight_1[235]), .B1(
        n17815), .Y(n17469) );
  AOI22XL U21599 ( .A0(weight_1[223]), .A1(n17811), .B0(weight_1[145]), .B1(
        n17822), .Y(n17468) );
  AOI22XL U21600 ( .A0(weight_1[379]), .A1(n17821), .B0(weight_1[355]), .B1(
        n17827), .Y(n17467) );
  NAND4XL U21601 ( .A(n17470), .B(n17469), .C(n17468), .D(n17467), .Y(n17471)
         );
  NOR4XL U21602 ( .A(n17474), .B(n17473), .C(n17472), .D(n17471), .Y(n17496)
         );
  AOI22XL U21603 ( .A0(n16744), .A1(weight_1[79]), .B0(weight_1[277]), .B1(
        n17802), .Y(n17478) );
  AOI22XL U21604 ( .A0(weight_1[271]), .A1(n17877), .B0(weight_1[241]), .B1(
        n17797), .Y(n17477) );
  AOI22XL U21605 ( .A0(n21762), .A1(weight_1[7]), .B0(weight_1[157]), .B1(
        n17863), .Y(n17476) );
  AOI22XL U21606 ( .A0(weight_1[295]), .A1(n17798), .B0(weight_1[199]), .B1(
        n17884), .Y(n17475) );
  NAND4XL U21607 ( .A(n17478), .B(n17477), .C(n17476), .D(n17475), .Y(n17494)
         );
  AOI22XL U21608 ( .A0(n26082), .A1(weight_1[319]), .B0(weight_1[91]), .B1(
        n17897), .Y(n17482) );
  AOI22XL U21609 ( .A0(n21748), .A1(weight_1[307]), .B0(weight_1[25]), .B1(
        n17873), .Y(n17481) );
  AOI22XL U21610 ( .A0(weight_1[139]), .A1(n17875), .B0(weight_1[55]), .B1(
        n17791), .Y(n17480) );
  AOI22XL U21611 ( .A0(n21766), .A1(weight_1[313]), .B0(weight_1[49]), .B1(
        n17789), .Y(n17479) );
  NAND4XL U21612 ( .A(n17482), .B(n17481), .C(n17480), .D(n17479), .Y(n17493)
         );
  AOI22XL U21613 ( .A0(weight_1[103]), .A1(n17887), .B0(weight_1[37]), .B1(
        n17874), .Y(n17486) );
  AOI22XL U21614 ( .A0(weight_1[121]), .A1(n17801), .B0(weight_1[73]), .B1(
        n17799), .Y(n17485) );
  AOI22XL U21615 ( .A0(weight_1[181]), .A1(n17790), .B0(weight_1[151]), .B1(
        n17868), .Y(n17484) );
  AOI22XL U21616 ( .A0(n21764), .A1(weight_1[13]), .B0(weight_1[163]), .B1(
        n17888), .Y(n17483) );
  NAND4XL U21617 ( .A(n17486), .B(n17485), .C(n17484), .D(n17483), .Y(n17492)
         );
  AOI22XL U21618 ( .A0(weight_1[385]), .A1(n17800), .B0(weight_1[61]), .B1(
        n17883), .Y(n17490) );
  AOI22XL U21619 ( .A0(weight_1[43]), .A1(n17803), .B0(weight_1[31]), .B1(
        n17867), .Y(n17489) );
  AOI22XL U21620 ( .A0(weight_1[301]), .A1(n17787), .B0(weight_1[247]), .B1(
        n17896), .Y(n17488) );
  AOI22XL U21621 ( .A0(weight_1[259]), .A1(n17788), .B0(weight_1[67]), .B1(
        n17865), .Y(n17487) );
  NAND4XL U21622 ( .A(n17490), .B(n17489), .C(n17488), .D(n17487), .Y(n17491)
         );
  NOR4XL U21623 ( .A(n17494), .B(n17493), .C(n17492), .D(n17491), .Y(n17495)
         );
  OAI2BB1XL U21624 ( .A0N(n17496), .A1N(n17495), .B0(n19182), .Y(n17497) );
  NAND4X1 U21625 ( .A(n17500), .B(n17499), .C(n17498), .D(n17497), .Y(n20629)
         );
  NAND2XL U21626 ( .A(n33554), .B(n20629), .Y(DP_OP_5167J1_123_9881_n56) );
  NAND2XL U21627 ( .A(n33553), .B(n20645), .Y(DP_OP_5167J1_123_9881_n76) );
  NAND2XL U21628 ( .A(n33554), .B(n20628), .Y(DP_OP_5167J1_123_9881_n55) );
  NAND2XL U21629 ( .A(n33554), .B(n17506), .Y(DP_OP_5167J1_123_9881_n54) );
  NAND2XL U21630 ( .A(n33553), .B(n17918), .Y(DP_OP_5167J1_123_9881_n58) );
  NAND2XL U21631 ( .A(n33554), .B(n17507), .Y(DP_OP_5167J1_123_9881_n53) );
  INVXL U21632 ( .A(affine_1[15]), .Y(DP_OP_5167J1_123_9881_n33) );
  AND2XL U21633 ( .A(n20629), .B(n20646), .Y(n17501) );
  AND2XL U21634 ( .A(n20629), .B(n17918), .Y(n17504) );
  AND2XL U21635 ( .A(n17506), .B(n20648), .Y(n17503) );
  ADDHXL U21636 ( .A(affine_1[13]), .B(n17501), .CO(n17502), .S(
        DP_OP_5167J1_123_9881_n45) );
  ADDFX1 U21637 ( .A(n17504), .B(n17503), .CI(n17502), .CO(
        DP_OP_5167J1_123_9881_n37), .S(DP_OP_5167J1_123_9881_n38) );
  AND2XL U21638 ( .A(n20645), .B(n17506), .Y(DP_OP_5167J1_123_9881_n78) );
  AND2XL U21639 ( .A(n20634), .B(n17918), .Y(DP_OP_5167J1_123_9881_n63) );
  AND2XL U21640 ( .A(n17506), .B(n20646), .Y(DP_OP_5167J1_123_9881_n66) );
  AND2XL U21641 ( .A(n17507), .B(n20648), .Y(DP_OP_5167J1_123_9881_n71) );
  AND2XL U21642 ( .A(n17507), .B(n17918), .Y(n17509) );
  NAND2XL U21643 ( .A(n33553), .B(n20646), .Y(n17508) );
  AOI22XL U21644 ( .A0(n21764), .A1(weight_1[10]), .B0(weight_1[382]), .B1(
        n17800), .Y(n17513) );
  AOI22XL U21645 ( .A0(weight_1[52]), .A1(n17791), .B0(weight_1[28]), .B1(
        n17867), .Y(n17512) );
  AOI22XL U21646 ( .A0(weight_1[274]), .A1(n17802), .B0(weight_1[130]), .B1(
        n17894), .Y(n17511) );
  AOI22XL U21647 ( .A0(weight_1[298]), .A1(n17787), .B0(weight_1[112]), .B1(
        n17792), .Y(n17510) );
  NAND4XL U21648 ( .A(n17513), .B(n17512), .C(n17511), .D(n17510), .Y(n17529)
         );
  AOI22XL U21649 ( .A0(weight_1[214]), .A1(n17878), .B0(weight_1[124]), .B1(
        n17895), .Y(n17517) );
  AOI22XL U21650 ( .A0(weight_1[268]), .A1(n17877), .B0(weight_1[154]), .B1(
        n17863), .Y(n17516) );
  AOI22XL U21651 ( .A0(weight_1[202]), .A1(n17898), .B0(weight_1[106]), .B1(
        n17876), .Y(n17515) );
  AOI22XL U21652 ( .A0(weight_1[208]), .A1(n17804), .B0(weight_1[184]), .B1(
        n17866), .Y(n17514) );
  NAND4XL U21653 ( .A(n17517), .B(n17516), .C(n17515), .D(n17514), .Y(n17528)
         );
  AOI22XL U21654 ( .A0(weight_1[370]), .A1(n17810), .B0(weight_1[232]), .B1(
        n17815), .Y(n17521) );
  AOI22XL U21655 ( .A0(weight_1[328]), .A1(n17814), .B0(weight_1[220]), .B1(
        n17811), .Y(n17520) );
  AOI22XL U21656 ( .A0(weight_1[346]), .A1(n17816), .B0(weight_1[334]), .B1(
        n17823), .Y(n17519) );
  AOI22XL U21657 ( .A0(weight_1[358]), .A1(n17825), .B0(weight_1[190]), .B1(
        n17813), .Y(n17518) );
  NAND4XL U21658 ( .A(n17521), .B(n17520), .C(n17519), .D(n17518), .Y(n17527)
         );
  AOI22XL U21659 ( .A0(weight_1[340]), .A1(n17812), .B0(weight_1[292]), .B1(
        n17798), .Y(n17525) );
  AOI22XL U21660 ( .A0(weight_1[226]), .A1(n17824), .B0(weight_1[142]), .B1(
        n17822), .Y(n17524) );
  AOI22XL U21661 ( .A0(weight_1[352]), .A1(n17827), .B0(weight_1[286]), .B1(
        n17826), .Y(n17523) );
  AOI22XL U21662 ( .A0(weight_1[376]), .A1(n17821), .B0(weight_1[364]), .B1(
        n17809), .Y(n17522) );
  NAND4XL U21663 ( .A(n17525), .B(n17524), .C(n17523), .D(n17522), .Y(n17526)
         );
  NOR4XL U21664 ( .A(n17529), .B(n17528), .C(n17527), .D(n17526), .Y(n17562)
         );
  INVXL U21665 ( .A(weight_1[424]), .Y(n32753) );
  INVXL U21666 ( .A(n17755), .Y(n17839) );
  OAI22XL U21667 ( .A0(n32760), .A1(n17749), .B0(n32753), .B1(n17839), .Y(
        n17539) );
  INVXL U21668 ( .A(weight_1[406]), .Y(n32382) );
  INVXL U21669 ( .A(n17840), .Y(n17583) );
  OAI22XL U21670 ( .A0(n32384), .A1(n17746), .B0(n32382), .B1(n17583), .Y(
        n17538) );
  INVXL U21671 ( .A(weight_1[466]), .Y(n32757) );
  AOI22XL U21672 ( .A0(weight_1[484]), .A1(n17841), .B0(weight_1[430]), .B1(
        n17752), .Y(n17531) );
  AOI22XL U21673 ( .A0(weight_1[478]), .A1(n17843), .B0(weight_1[460]), .B1(
        n17691), .Y(n17530) );
  OAI211XL U21674 ( .A0(n32757), .A1(n17694), .B0(n17531), .C0(n17530), .Y(
        n17537) );
  AOI22XL U21675 ( .A0(weight_1[454]), .A1(n17852), .B0(weight_1[436]), .B1(
        n17848), .Y(n17535) );
  AOI22XL U21676 ( .A0(weight_1[448]), .A1(n17753), .B0(weight_1[388]), .B1(
        n17754), .Y(n17534) );
  AOI22XL U21677 ( .A0(weight_1[412]), .A1(n17854), .B0(weight_1[400]), .B1(
        n17851), .Y(n17533) );
  AOI22XL U21678 ( .A0(weight_1[418]), .A1(n17847), .B0(weight_1[394]), .B1(
        n17853), .Y(n17532) );
  NAND4XL U21679 ( .A(n17535), .B(n17534), .C(n17533), .D(n17532), .Y(n17536)
         );
  NOR4XL U21680 ( .A(n17539), .B(n17538), .C(n17537), .D(n17536), .Y(n17561)
         );
  AOI22XL U21681 ( .A0(weight_1[64]), .A1(n17865), .B0(weight_1[22]), .B1(
        n17873), .Y(n17543) );
  AOI22XL U21682 ( .A0(weight_1[178]), .A1(n17790), .B0(weight_1[88]), .B1(
        n17897), .Y(n17542) );
  AOI22XL U21683 ( .A0(weight_1[244]), .A1(n17896), .B0(weight_1[172]), .B1(
        n16724), .Y(n17541) );
  AOI22XL U21684 ( .A0(weight_1[256]), .A1(n17788), .B0(weight_1[70]), .B1(
        n17799), .Y(n17540) );
  NAND4XL U21685 ( .A(n17543), .B(n17542), .C(n17541), .D(n17540), .Y(n17559)
         );
  AOI22XL U21686 ( .A0(weight_1[148]), .A1(n17868), .B0(weight_1[100]), .B1(
        n17887), .Y(n17547) );
  AOI22XL U21687 ( .A0(weight_1[250]), .A1(n17886), .B0(weight_1[160]), .B1(
        n17888), .Y(n17546) );
  AOI22XL U21688 ( .A0(weight_1[196]), .A1(n17884), .B0(weight_1[16]), .B1(
        n17893), .Y(n17545) );
  AOI22XL U21689 ( .A0(n21762), .A1(weight_1[4]), .B0(weight_1[58]), .B1(
        n17883), .Y(n17544) );
  NAND4XL U21690 ( .A(n17547), .B(n17546), .C(n17545), .D(n17544), .Y(n17558)
         );
  AOI22XL U21691 ( .A0(n26059), .A1(weight_1[322]), .B0(weight_1[136]), .B1(
        n17875), .Y(n17551) );
  AOI22XL U21692 ( .A0(weight_1[118]), .A1(n17801), .B0(weight_1[34]), .B1(
        n17874), .Y(n17550) );
  AOI22XL U21693 ( .A0(weight_1[166]), .A1(n17899), .B0(weight_1[46]), .B1(
        n17789), .Y(n17549) );
  AOI22XL U21694 ( .A0(n21748), .A1(weight_1[304]), .B0(weight_1[40]), .B1(
        n17803), .Y(n17548) );
  NAND4XL U21695 ( .A(n17551), .B(n17550), .C(n17549), .D(n17548), .Y(n17557)
         );
  AOI22XL U21696 ( .A0(n16744), .A1(weight_1[76]), .B0(n21766), .B1(
        weight_1[310]), .Y(n17555) );
  AOI22XL U21697 ( .A0(weight_1[280]), .A1(n17900), .B0(weight_1[94]), .B1(
        n17885), .Y(n17554) );
  AOI22XL U21698 ( .A0(weight_1[262]), .A1(n17864), .B0(weight_1[238]), .B1(
        n17797), .Y(n17553) );
  AOI22XL U21699 ( .A0(n26082), .A1(weight_1[316]), .B0(n21999), .B1(
        weight_1[82]), .Y(n17552) );
  NAND4XL U21700 ( .A(n17555), .B(n17554), .C(n17553), .D(n17552), .Y(n17556)
         );
  NOR4XL U21701 ( .A(n17559), .B(n17558), .C(n17557), .D(n17556), .Y(n17560)
         );
  AOI32XL U21702 ( .A0(n17562), .A1(n17561), .A2(n17560), .B0(cursor[6]), .B1(
        n17561), .Y(n17919) );
  NAND2XL U21703 ( .A(n20645), .B(n17919), .Y(n17917) );
  NAND2BXL U21704 ( .AN(affine_1[4]), .B(n17917), .Y(DP_OP_5168J1_124_9881_n39) );
  AOI22XL U21705 ( .A0(weight_1[183]), .A1(n17866), .B0(weight_1[117]), .B1(
        n17801), .Y(n17566) );
  AOI22XL U21706 ( .A0(weight_1[57]), .A1(n17883), .B0(weight_1[33]), .B1(
        n17874), .Y(n17565) );
  AOI22XL U21707 ( .A0(weight_1[123]), .A1(n17895), .B0(weight_1[69]), .B1(
        n17799), .Y(n17564) );
  AOI22XL U21708 ( .A0(n21766), .A1(weight_1[309]), .B0(weight_1[21]), .B1(
        n17873), .Y(n17563) );
  NAND4XL U21709 ( .A(n17566), .B(n17565), .C(n17564), .D(n17563), .Y(n17582)
         );
  AOI22XL U21710 ( .A0(n21762), .A1(weight_1[3]), .B0(weight_1[129]), .B1(
        n17894), .Y(n17570) );
  AOI22XL U21711 ( .A0(weight_1[153]), .A1(n17863), .B0(weight_1[99]), .B1(
        n17887), .Y(n17569) );
  AOI22XL U21712 ( .A0(weight_1[291]), .A1(n17798), .B0(weight_1[15]), .B1(
        n17893), .Y(n17568) );
  AOI22XL U21713 ( .A0(n26082), .A1(weight_1[315]), .B0(weight_1[105]), .B1(
        n17876), .Y(n17567) );
  NAND4XL U21714 ( .A(n17570), .B(n17569), .C(n17568), .D(n17567), .Y(n17581)
         );
  AOI22XL U21715 ( .A0(weight_1[351]), .A1(n17827), .B0(weight_1[345]), .B1(
        n17816), .Y(n17574) );
  AOI22XL U21716 ( .A0(weight_1[369]), .A1(n17810), .B0(weight_1[141]), .B1(
        n17822), .Y(n17573) );
  AOI22XL U21717 ( .A0(weight_1[357]), .A1(n17825), .B0(weight_1[189]), .B1(
        n17813), .Y(n17572) );
  AOI22XL U21718 ( .A0(weight_1[285]), .A1(n17826), .B0(weight_1[225]), .B1(
        n17824), .Y(n17571) );
  NAND4XL U21719 ( .A(n17574), .B(n17573), .C(n17572), .D(n17571), .Y(n17580)
         );
  AOI22XL U21720 ( .A0(weight_1[327]), .A1(n17814), .B0(weight_1[39]), .B1(
        n17803), .Y(n17578) );
  AOI22XL U21721 ( .A0(weight_1[375]), .A1(n17821), .B0(weight_1[363]), .B1(
        n17809), .Y(n17577) );
  AOI22XL U21722 ( .A0(weight_1[339]), .A1(n17812), .B0(weight_1[333]), .B1(
        n17823), .Y(n17576) );
  AOI22XL U21723 ( .A0(weight_1[231]), .A1(n17815), .B0(weight_1[219]), .B1(
        n17811), .Y(n17575) );
  NAND4XL U21724 ( .A(n17578), .B(n17577), .C(n17576), .D(n17575), .Y(n17579)
         );
  NOR4XL U21725 ( .A(n17582), .B(n17581), .C(n17580), .D(n17579), .Y(n17616)
         );
  INVXL U21726 ( .A(weight_1[435]), .Y(n32499) );
  INVXL U21727 ( .A(weight_1[399]), .Y(n32510) );
  OAI22XL U21728 ( .A0(n32499), .A1(n17690), .B0(n32510), .B1(n17748), .Y(
        n17593) );
  INVXL U21729 ( .A(weight_1[405]), .Y(n32509) );
  OAI22XL U21730 ( .A0(n32484), .A1(n17837), .B0(n32509), .B1(n17583), .Y(
        n17592) );
  AOI22XL U21731 ( .A0(weight_1[483]), .A1(n17841), .B0(weight_1[423]), .B1(
        n17755), .Y(n17585) );
  AOI22XL U21732 ( .A0(weight_1[477]), .A1(n17843), .B0(weight_1[459]), .B1(
        n17691), .Y(n17584) );
  OAI211XL U21733 ( .A0(n32473), .A1(n17694), .B0(n17585), .C0(n17584), .Y(
        n17591) );
  AOI22XL U21734 ( .A0(weight_1[471]), .A1(n17850), .B0(weight_1[393]), .B1(
        n17853), .Y(n17589) );
  AOI22XL U21735 ( .A0(weight_1[453]), .A1(n17852), .B0(weight_1[387]), .B1(
        n17754), .Y(n17588) );
  AOI22XL U21736 ( .A0(weight_1[429]), .A1(n17752), .B0(weight_1[411]), .B1(
        n17854), .Y(n17587) );
  AOI22XL U21737 ( .A0(weight_1[441]), .A1(n17849), .B0(weight_1[417]), .B1(
        n17847), .Y(n17586) );
  NAND4XL U21738 ( .A(n17589), .B(n17588), .C(n17587), .D(n17586), .Y(n17590)
         );
  NOR4XL U21739 ( .A(n17593), .B(n17592), .C(n17591), .D(n17590), .Y(n17615)
         );
  AOI22XL U21740 ( .A0(weight_1[261]), .A1(n17864), .B0(weight_1[249]), .B1(
        n17886), .Y(n17597) );
  AOI22XL U21741 ( .A0(weight_1[279]), .A1(n17900), .B0(weight_1[171]), .B1(
        n16724), .Y(n17596) );
  AOI22XL U21742 ( .A0(n26059), .A1(weight_1[321]), .B0(weight_1[267]), .B1(
        n17877), .Y(n17595) );
  AOI22XL U21743 ( .A0(weight_1[243]), .A1(n17896), .B0(weight_1[51]), .B1(
        n17791), .Y(n17594) );
  NAND4XL U21744 ( .A(n17597), .B(n17596), .C(n17595), .D(n17594), .Y(n17613)
         );
  AOI22XL U21745 ( .A0(n21748), .A1(weight_1[303]), .B0(weight_1[111]), .B1(
        n17792), .Y(n17601) );
  AOI22XL U21746 ( .A0(weight_1[237]), .A1(n17797), .B0(weight_1[147]), .B1(
        n17868), .Y(n17600) );
  AOI22XL U21747 ( .A0(n21764), .A1(weight_1[9]), .B0(weight_1[45]), .B1(
        n17789), .Y(n17599) );
  AOI22XL U21748 ( .A0(weight_1[201]), .A1(n17898), .B0(weight_1[93]), .B1(
        n17885), .Y(n17598) );
  NAND4XL U21749 ( .A(n17601), .B(n17600), .C(n17599), .D(n17598), .Y(n17612)
         );
  AOI22XL U21750 ( .A0(weight_1[255]), .A1(n17788), .B0(weight_1[213]), .B1(
        n17878), .Y(n17605) );
  AOI22XL U21751 ( .A0(weight_1[195]), .A1(n17884), .B0(weight_1[135]), .B1(
        n17875), .Y(n17604) );
  AOI22XL U21752 ( .A0(n21999), .A1(weight_1[81]), .B0(weight_1[273]), .B1(
        n17802), .Y(n17603) );
  AOI22XL U21753 ( .A0(weight_1[63]), .A1(n17865), .B0(weight_1[27]), .B1(
        n17867), .Y(n17602) );
  NAND4XL U21754 ( .A(n17605), .B(n17604), .C(n17603), .D(n17602), .Y(n17611)
         );
  AOI22XL U21755 ( .A0(weight_1[381]), .A1(n17800), .B0(weight_1[87]), .B1(
        n17897), .Y(n17609) );
  AOI22XL U21756 ( .A0(weight_1[297]), .A1(n17787), .B0(weight_1[165]), .B1(
        n17899), .Y(n17608) );
  AOI22XL U21757 ( .A0(n16744), .A1(weight_1[75]), .B0(weight_1[159]), .B1(
        n17888), .Y(n17607) );
  AOI22XL U21758 ( .A0(weight_1[207]), .A1(n17804), .B0(weight_1[177]), .B1(
        n17790), .Y(n17606) );
  NAND4XL U21759 ( .A(n17609), .B(n17608), .C(n17607), .D(n17606), .Y(n17610)
         );
  NOR4XL U21760 ( .A(n17613), .B(n17612), .C(n17611), .D(n17610), .Y(n17614)
         );
  AND2XL U21761 ( .A(n17916), .B(n17918), .Y(DP_OP_5168J1_124_9881_n60) );
  AOI22XL U21762 ( .A0(weight_1[152]), .A1(n17863), .B0(weight_1[92]), .B1(
        n17885), .Y(n17620) );
  AOI22XL U21763 ( .A0(n21748), .A1(weight_1[302]), .B0(weight_1[56]), .B1(
        n17883), .Y(n17619) );
  AOI22XL U21764 ( .A0(weight_1[62]), .A1(n17865), .B0(weight_1[38]), .B1(
        n17803), .Y(n17618) );
  AOI22XL U21765 ( .A0(weight_1[266]), .A1(n17877), .B0(weight_1[14]), .B1(
        n17893), .Y(n17617) );
  NAND4XL U21766 ( .A(n17620), .B(n17619), .C(n17618), .D(n17617), .Y(n17636)
         );
  AOI22XL U21767 ( .A0(n26082), .A1(weight_1[314]), .B0(n21999), .B1(
        weight_1[80]), .Y(n17624) );
  AOI22XL U21768 ( .A0(weight_1[110]), .A1(n17792), .B0(weight_1[86]), .B1(
        n17897), .Y(n17623) );
  AOI22XL U21769 ( .A0(weight_1[158]), .A1(n17888), .B0(weight_1[26]), .B1(
        n17867), .Y(n17622) );
  AOI22XL U21770 ( .A0(weight_1[296]), .A1(n17787), .B0(weight_1[44]), .B1(
        n17789), .Y(n17621) );
  NAND4XL U21771 ( .A(n17624), .B(n17623), .C(n17622), .D(n17621), .Y(n17635)
         );
  AOI22XL U21772 ( .A0(weight_1[374]), .A1(n17821), .B0(weight_1[224]), .B1(
        n17824), .Y(n17628) );
  AOI22XL U21773 ( .A0(weight_1[284]), .A1(n17826), .B0(weight_1[188]), .B1(
        n17813), .Y(n17627) );
  AOI22XL U21774 ( .A0(weight_1[368]), .A1(n17810), .B0(weight_1[326]), .B1(
        n17814), .Y(n17626) );
  AOI22XL U21775 ( .A0(weight_1[332]), .A1(n17823), .B0(weight_1[218]), .B1(
        n17811), .Y(n17625) );
  NAND4XL U21776 ( .A(n17628), .B(n17627), .C(n17626), .D(n17625), .Y(n17634)
         );
  AOI22XL U21777 ( .A0(n21762), .A1(weight_1[2]), .B0(weight_1[230]), .B1(
        n17815), .Y(n17632) );
  AOI22XL U21778 ( .A0(weight_1[356]), .A1(n17825), .B0(weight_1[140]), .B1(
        n17822), .Y(n17631) );
  AOI22XL U21779 ( .A0(weight_1[362]), .A1(n17809), .B0(weight_1[350]), .B1(
        n17827), .Y(n17630) );
  AOI22XL U21780 ( .A0(weight_1[344]), .A1(n17816), .B0(weight_1[338]), .B1(
        n17812), .Y(n17629) );
  NAND4XL U21781 ( .A(n17632), .B(n17631), .C(n17630), .D(n17629), .Y(n17633)
         );
  NOR4XL U21782 ( .A(n17636), .B(n17635), .C(n17634), .D(n17633), .Y(n17669)
         );
  INVXL U21783 ( .A(weight_1[386]), .Y(n32398) );
  OAI2BB2XL U21784 ( .B0(n32398), .B1(n17838), .A0N(weight_1[410]), .A1N(
        n17854), .Y(n17646) );
  INVXL U21785 ( .A(weight_1[428]), .Y(n32390) );
  INVXL U21786 ( .A(n17752), .Y(n17836) );
  OAI22XL U21787 ( .A0(n32379), .A1(n17747), .B0(n32390), .B1(n17836), .Y(
        n17645) );
  INVXL U21788 ( .A(weight_1[458]), .Y(n32372) );
  AOI22XL U21789 ( .A0(weight_1[482]), .A1(n17841), .B0(weight_1[416]), .B1(
        n17847), .Y(n17638) );
  AOI22XL U21790 ( .A0(weight_1[476]), .A1(n17843), .B0(weight_1[464]), .B1(
        n17842), .Y(n17637) );
  OAI211XL U21791 ( .A0(n32372), .A1(n17846), .B0(n17638), .C0(n17637), .Y(
        n17644) );
  AOI22XL U21792 ( .A0(weight_1[446]), .A1(n17753), .B0(weight_1[440]), .B1(
        n17849), .Y(n17642) );
  AOI22XL U21793 ( .A0(weight_1[434]), .A1(n17848), .B0(weight_1[398]), .B1(
        n17851), .Y(n17641) );
  AOI22XL U21794 ( .A0(weight_1[422]), .A1(n17755), .B0(weight_1[392]), .B1(
        n17853), .Y(n17640) );
  AOI22XL U21795 ( .A0(weight_1[470]), .A1(n17850), .B0(weight_1[404]), .B1(
        n17840), .Y(n17639) );
  NAND4XL U21796 ( .A(n17642), .B(n17641), .C(n17640), .D(n17639), .Y(n17643)
         );
  NOR4XL U21797 ( .A(n17646), .B(n17645), .C(n17644), .D(n17643), .Y(n17668)
         );
  AOI22XL U21798 ( .A0(n26059), .A1(weight_1[320]), .B0(weight_1[104]), .B1(
        n17876), .Y(n17650) );
  AOI22XL U21799 ( .A0(n21766), .A1(weight_1[308]), .B0(weight_1[164]), .B1(
        n17899), .Y(n17649) );
  AOI22XL U21800 ( .A0(weight_1[242]), .A1(n17896), .B0(weight_1[236]), .B1(
        n17797), .Y(n17648) );
  AOI22XL U21801 ( .A0(weight_1[32]), .A1(n17874), .B0(weight_1[20]), .B1(
        n17873), .Y(n17647) );
  NAND4XL U21802 ( .A(n17650), .B(n17649), .C(n17648), .D(n17647), .Y(n17666)
         );
  AOI22XL U21803 ( .A0(weight_1[260]), .A1(n17864), .B0(weight_1[116]), .B1(
        n17801), .Y(n17654) );
  AOI22XL U21804 ( .A0(weight_1[146]), .A1(n17868), .B0(weight_1[50]), .B1(
        n17791), .Y(n17653) );
  AOI22XL U21805 ( .A0(weight_1[212]), .A1(n17878), .B0(weight_1[200]), .B1(
        n17898), .Y(n17652) );
  AOI22XL U21806 ( .A0(weight_1[380]), .A1(n17800), .B0(weight_1[170]), .B1(
        n16724), .Y(n17651) );
  NAND4XL U21807 ( .A(n17654), .B(n17653), .C(n17652), .D(n17651), .Y(n17665)
         );
  AOI22XL U21808 ( .A0(weight_1[254]), .A1(n17788), .B0(weight_1[98]), .B1(
        n17887), .Y(n17658) );
  AOI22XL U21809 ( .A0(weight_1[248]), .A1(n17886), .B0(weight_1[182]), .B1(
        n17866), .Y(n17657) );
  AOI22XL U21810 ( .A0(weight_1[278]), .A1(n17900), .B0(weight_1[194]), .B1(
        n17884), .Y(n17656) );
  AOI22XL U21811 ( .A0(n21764), .A1(weight_1[8]), .B0(weight_1[128]), .B1(
        n17894), .Y(n17655) );
  NAND4XL U21812 ( .A(n17658), .B(n17657), .C(n17656), .D(n17655), .Y(n17664)
         );
  AOI22XL U21813 ( .A0(weight_1[272]), .A1(n17802), .B0(weight_1[68]), .B1(
        n17799), .Y(n17662) );
  AOI22XL U21814 ( .A0(weight_1[176]), .A1(n17790), .B0(weight_1[134]), .B1(
        n17875), .Y(n17661) );
  AOI22XL U21815 ( .A0(n16744), .A1(weight_1[74]), .B0(weight_1[206]), .B1(
        n17804), .Y(n17660) );
  AOI22XL U21816 ( .A0(weight_1[290]), .A1(n17798), .B0(weight_1[122]), .B1(
        n17895), .Y(n17659) );
  NAND4XL U21817 ( .A(n17662), .B(n17661), .C(n17660), .D(n17659), .Y(n17663)
         );
  NOR4XL U21818 ( .A(n17666), .B(n17665), .C(n17664), .D(n17663), .Y(n17667)
         );
  AND2XL U21819 ( .A(n20644), .B(n17918), .Y(DP_OP_5168J1_124_9881_n61) );
  AND2XL U21820 ( .A(n20644), .B(n20646), .Y(DP_OP_5168J1_124_9881_n67) );
  AND2XL U21821 ( .A(n20644), .B(n20648), .Y(DP_OP_5168J1_124_9881_n73) );
  AOI22XL U21822 ( .A0(weight_1[203]), .A1(n17898), .B0(weight_1[35]), .B1(
        n17874), .Y(n17673) );
  AOI22XL U21823 ( .A0(weight_1[155]), .A1(n17863), .B0(weight_1[59]), .B1(
        n17883), .Y(n17672) );
  AOI22XL U21824 ( .A0(weight_1[281]), .A1(n17900), .B0(weight_1[275]), .B1(
        n17802), .Y(n17671) );
  AOI22XL U21825 ( .A0(weight_1[29]), .A1(n17867), .B0(weight_1[17]), .B1(
        n17893), .Y(n17670) );
  NAND4XL U21826 ( .A(n17673), .B(n17672), .C(n17671), .D(n17670), .Y(n17689)
         );
  AOI22XL U21827 ( .A0(n21762), .A1(weight_1[5]), .B0(n21766), .B1(
        weight_1[311]), .Y(n17677) );
  AOI22XL U21828 ( .A0(weight_1[179]), .A1(n17790), .B0(weight_1[89]), .B1(
        n17897), .Y(n17676) );
  AOI22XL U21829 ( .A0(weight_1[209]), .A1(n17804), .B0(weight_1[41]), .B1(
        n17803), .Y(n17675) );
  AOI22XL U21830 ( .A0(weight_1[269]), .A1(n17877), .B0(weight_1[257]), .B1(
        n17788), .Y(n17674) );
  NAND4XL U21831 ( .A(n17677), .B(n17676), .C(n17675), .D(n17674), .Y(n17688)
         );
  AOI22XL U21832 ( .A0(weight_1[233]), .A1(n17815), .B0(weight_1[221]), .B1(
        n17811), .Y(n17681) );
  AOI22XL U21833 ( .A0(weight_1[365]), .A1(n17809), .B0(weight_1[287]), .B1(
        n17826), .Y(n17680) );
  AOI22XL U21834 ( .A0(weight_1[371]), .A1(n17810), .B0(weight_1[329]), .B1(
        n17814), .Y(n17679) );
  AOI22XL U21835 ( .A0(weight_1[353]), .A1(n17827), .B0(weight_1[347]), .B1(
        n17816), .Y(n17678) );
  NAND4XL U21836 ( .A(n17681), .B(n17680), .C(n17679), .D(n17678), .Y(n17687)
         );
  AOI22XL U21837 ( .A0(weight_1[377]), .A1(n17821), .B0(weight_1[161]), .B1(
        n17888), .Y(n17685) );
  AOI22XL U21838 ( .A0(weight_1[341]), .A1(n17812), .B0(weight_1[191]), .B1(
        n17813), .Y(n17684) );
  AOI22XL U21839 ( .A0(weight_1[335]), .A1(n17823), .B0(weight_1[143]), .B1(
        n17822), .Y(n17683) );
  AOI22XL U21840 ( .A0(weight_1[359]), .A1(n17825), .B0(weight_1[227]), .B1(
        n17824), .Y(n17682) );
  NAND4XL U21841 ( .A(n17685), .B(n17684), .C(n17683), .D(n17682), .Y(n17686)
         );
  NOR4XL U21842 ( .A(n17689), .B(n17688), .C(n17687), .D(n17686), .Y(n17725)
         );
  INVXL U21843 ( .A(weight_1[437]), .Y(n32921) );
  OAI2BB2XL U21844 ( .B0(n32921), .B1(n17690), .A0N(weight_1[419]), .A1N(
        n17847), .Y(n17702) );
  INVXL U21845 ( .A(weight_1[473]), .Y(n32905) );
  INVXL U21846 ( .A(weight_1[443]), .Y(n32923) );
  OAI22XL U21847 ( .A0(n32905), .A1(n17749), .B0(n32923), .B1(n17746), .Y(
        n17701) );
  AOI22XL U21848 ( .A0(weight_1[485]), .A1(n17841), .B0(weight_1[395]), .B1(
        n17853), .Y(n17693) );
  AOI22XL U21849 ( .A0(weight_1[479]), .A1(n17843), .B0(weight_1[461]), .B1(
        n17691), .Y(n17692) );
  OAI211XL U21850 ( .A0(n32906), .A1(n17694), .B0(n17693), .C0(n17692), .Y(
        n17700) );
  AOI22XL U21851 ( .A0(weight_1[455]), .A1(n17852), .B0(weight_1[413]), .B1(
        n17854), .Y(n17698) );
  AOI22XL U21852 ( .A0(weight_1[449]), .A1(n17753), .B0(weight_1[431]), .B1(
        n17752), .Y(n17697) );
  AOI22XL U21853 ( .A0(weight_1[407]), .A1(n17840), .B0(weight_1[389]), .B1(
        n17754), .Y(n17696) );
  AOI22XL U21854 ( .A0(weight_1[425]), .A1(n17755), .B0(weight_1[401]), .B1(
        n17851), .Y(n17695) );
  NAND4XL U21855 ( .A(n17698), .B(n17697), .C(n17696), .D(n17695), .Y(n17699)
         );
  NOR4XL U21856 ( .A(n17702), .B(n17701), .C(n17700), .D(n17699), .Y(n17724)
         );
  AOI22XL U21857 ( .A0(weight_1[185]), .A1(n17866), .B0(weight_1[53]), .B1(
        n17791), .Y(n17706) );
  AOI22XL U21858 ( .A0(weight_1[251]), .A1(n17886), .B0(weight_1[95]), .B1(
        n17885), .Y(n17705) );
  AOI22XL U21859 ( .A0(weight_1[167]), .A1(n17899), .B0(weight_1[125]), .B1(
        n17895), .Y(n17704) );
  AOI22XL U21860 ( .A0(weight_1[263]), .A1(n17864), .B0(weight_1[197]), .B1(
        n17884), .Y(n17703) );
  NAND4XL U21861 ( .A(n17706), .B(n17705), .C(n17704), .D(n17703), .Y(n17722)
         );
  AOI22XL U21862 ( .A0(n26059), .A1(weight_1[323]), .B0(n16744), .B1(
        weight_1[77]), .Y(n17710) );
  AOI22XL U21863 ( .A0(n21748), .A1(weight_1[305]), .B0(weight_1[299]), .B1(
        n17787), .Y(n17709) );
  AOI22XL U21864 ( .A0(weight_1[383]), .A1(n17800), .B0(weight_1[119]), .B1(
        n17801), .Y(n17708) );
  AOI22XL U21865 ( .A0(weight_1[137]), .A1(n17875), .B0(weight_1[23]), .B1(
        n17873), .Y(n17707) );
  NAND4XL U21866 ( .A(n17710), .B(n17709), .C(n17708), .D(n17707), .Y(n17721)
         );
  AOI22XL U21867 ( .A0(n21764), .A1(weight_1[11]), .B0(weight_1[173]), .B1(
        n16724), .Y(n17714) );
  AOI22XL U21868 ( .A0(weight_1[131]), .A1(n17894), .B0(weight_1[101]), .B1(
        n17887), .Y(n17713) );
  AOI22XL U21869 ( .A0(n21999), .A1(weight_1[83]), .B0(weight_1[65]), .B1(
        n17865), .Y(n17712) );
  AOI22XL U21870 ( .A0(weight_1[293]), .A1(n17798), .B0(weight_1[149]), .B1(
        n17868), .Y(n17711) );
  NAND4XL U21871 ( .A(n17714), .B(n17713), .C(n17712), .D(n17711), .Y(n17720)
         );
  AOI22XL U21872 ( .A0(weight_1[245]), .A1(n17896), .B0(weight_1[71]), .B1(
        n17799), .Y(n17718) );
  AOI22XL U21873 ( .A0(weight_1[239]), .A1(n17797), .B0(weight_1[113]), .B1(
        n17792), .Y(n17717) );
  AOI22XL U21874 ( .A0(weight_1[215]), .A1(n17878), .B0(weight_1[107]), .B1(
        n17876), .Y(n17716) );
  AOI22XL U21875 ( .A0(n26082), .A1(weight_1[317]), .B0(weight_1[47]), .B1(
        n17789), .Y(n17715) );
  NAND4XL U21876 ( .A(n17718), .B(n17717), .C(n17716), .D(n17715), .Y(n17719)
         );
  NOR4XL U21877 ( .A(n17722), .B(n17721), .C(n17720), .D(n17719), .Y(n17723)
         );
  AOI32XL U21878 ( .A0(n17725), .A1(n17724), .A2(n17723), .B0(cursor[6]), .B1(
        n17724), .Y(n33068) );
  NAND2XL U21879 ( .A(n33068), .B(n20648), .Y(DP_OP_5168J1_124_9881_n70) );
  AOI22XL U21880 ( .A0(n21766), .A1(weight_1[306]), .B0(weight_1[150]), .B1(
        n17863), .Y(n17729) );
  AOI22XL U21881 ( .A0(weight_1[234]), .A1(n17797), .B0(weight_1[18]), .B1(
        n17873), .Y(n17728) );
  AOI22XL U21882 ( .A0(weight_1[246]), .A1(n17886), .B0(weight_1[174]), .B1(
        n17790), .Y(n17727) );
  AOI22XL U21883 ( .A0(weight_1[264]), .A1(n17877), .B0(weight_1[90]), .B1(
        n17885), .Y(n17726) );
  NAND4XL U21884 ( .A(n17729), .B(n17728), .C(n17727), .D(n17726), .Y(n17745)
         );
  AOI22XL U21885 ( .A0(weight_1[204]), .A1(n17804), .B0(weight_1[180]), .B1(
        n17866), .Y(n17733) );
  AOI22XL U21886 ( .A0(weight_1[126]), .A1(n17894), .B0(weight_1[114]), .B1(
        n17801), .Y(n17732) );
  AOI22XL U21887 ( .A0(n16744), .A1(weight_1[72]), .B0(weight_1[168]), .B1(
        n16724), .Y(n17731) );
  AOI22XL U21888 ( .A0(weight_1[84]), .A1(n17897), .B0(weight_1[30]), .B1(
        n17874), .Y(n17730) );
  NAND4XL U21889 ( .A(n17733), .B(n17732), .C(n17731), .D(n17730), .Y(n17744)
         );
  AOI22XL U21890 ( .A0(weight_1[360]), .A1(n17809), .B0(weight_1[348]), .B1(
        n17827), .Y(n17737) );
  AOI22XL U21891 ( .A0(weight_1[366]), .A1(n17810), .B0(weight_1[222]), .B1(
        n17824), .Y(n17736) );
  AOI22XL U21892 ( .A0(weight_1[372]), .A1(n17821), .B0(weight_1[186]), .B1(
        n17813), .Y(n17735) );
  AOI22XL U21893 ( .A0(weight_1[342]), .A1(n17816), .B0(weight_1[216]), .B1(
        n17811), .Y(n17734) );
  NAND4XL U21894 ( .A(n17737), .B(n17736), .C(n17735), .D(n17734), .Y(n17743)
         );
  AOI22XL U21895 ( .A0(weight_1[330]), .A1(n17823), .B0(weight_1[66]), .B1(
        n17799), .Y(n17741) );
  AOI22XL U21896 ( .A0(weight_1[354]), .A1(n17825), .B0(weight_1[138]), .B1(
        n17822), .Y(n17740) );
  AOI22XL U21897 ( .A0(weight_1[282]), .A1(n17826), .B0(weight_1[228]), .B1(
        n17815), .Y(n17739) );
  AOI22XL U21898 ( .A0(weight_1[336]), .A1(n17812), .B0(weight_1[324]), .B1(
        n17814), .Y(n17738) );
  NAND4XL U21899 ( .A(n17741), .B(n17740), .C(n17739), .D(n17738), .Y(n17742)
         );
  NOR4XL U21900 ( .A(n17745), .B(n17744), .C(n17743), .D(n17742), .Y(n17786)
         );
  OAI22XL U21901 ( .A0(n26867), .A1(n17747), .B0(n26885), .B1(n17746), .Y(
        n17763) );
  OAI22XL U21902 ( .A0(n26907), .A1(n17749), .B0(n26912), .B1(n17748), .Y(
        n17762) );
  INVXL U21903 ( .A(weight_1[456]), .Y(n26880) );
  AOI22XL U21904 ( .A0(weight_1[480]), .A1(n17841), .B0(weight_1[432]), .B1(
        n17848), .Y(n17751) );
  AOI22XL U21905 ( .A0(weight_1[474]), .A1(n17843), .B0(weight_1[462]), .B1(
        n17842), .Y(n17750) );
  OAI211XL U21906 ( .A0(n26880), .A1(n17846), .B0(n17751), .C0(n17750), .Y(
        n17761) );
  AOI22XL U21907 ( .A0(weight_1[408]), .A1(n17854), .B0(weight_1[402]), .B1(
        n17840), .Y(n17759) );
  AOI22XL U21908 ( .A0(weight_1[444]), .A1(n17753), .B0(weight_1[426]), .B1(
        n17752), .Y(n17758) );
  AOI22XL U21909 ( .A0(weight_1[414]), .A1(n17847), .B0(weight_1[390]), .B1(
        n17853), .Y(n17757) );
  AOI22XL U21910 ( .A0(weight_1[420]), .A1(n17755), .B0(weight_1[384]), .B1(
        n17754), .Y(n17756) );
  NAND4XL U21911 ( .A(n17759), .B(n17758), .C(n17757), .D(n17756), .Y(n17760)
         );
  NOR4XL U21912 ( .A(n17763), .B(n17762), .C(n17761), .D(n17760), .Y(n17785)
         );
  AOI22XL U21913 ( .A0(n21764), .A1(weight_1[6]), .B0(weight_1[240]), .B1(
        n17896), .Y(n17767) );
  AOI22XL U21914 ( .A0(n21762), .A1(weight_1[0]), .B0(weight_1[198]), .B1(
        n17898), .Y(n17766) );
  AOI22XL U21915 ( .A0(weight_1[252]), .A1(n17788), .B0(weight_1[36]), .B1(
        n17803), .Y(n17765) );
  AOI22XL U21916 ( .A0(weight_1[60]), .A1(n17865), .B0(weight_1[54]), .B1(
        n17883), .Y(n17764) );
  NAND4XL U21917 ( .A(n17767), .B(n17766), .C(n17765), .D(n17764), .Y(n17783)
         );
  AOI22XL U21918 ( .A0(weight_1[258]), .A1(n17864), .B0(weight_1[156]), .B1(
        n17888), .Y(n17771) );
  AOI22XL U21919 ( .A0(n26059), .A1(weight_1[318]), .B0(weight_1[378]), .B1(
        n17800), .Y(n17770) );
  AOI22XL U21920 ( .A0(weight_1[132]), .A1(n17875), .B0(weight_1[96]), .B1(
        n17887), .Y(n17769) );
  AOI22XL U21921 ( .A0(weight_1[288]), .A1(n17798), .B0(weight_1[210]), .B1(
        n17878), .Y(n17768) );
  NAND4XL U21922 ( .A(n17771), .B(n17770), .C(n17769), .D(n17768), .Y(n17782)
         );
  AOI22XL U21923 ( .A0(n26082), .A1(weight_1[312]), .B0(weight_1[24]), .B1(
        n17867), .Y(n17775) );
  AOI22XL U21924 ( .A0(weight_1[276]), .A1(n17900), .B0(weight_1[162]), .B1(
        n17899), .Y(n17774) );
  AOI22XL U21925 ( .A0(n21748), .A1(weight_1[300]), .B0(weight_1[102]), .B1(
        n17876), .Y(n17773) );
  AOI22XL U21926 ( .A0(n21999), .A1(weight_1[78]), .B0(weight_1[48]), .B1(
        n17791), .Y(n17772) );
  NAND4XL U21927 ( .A(n17775), .B(n17774), .C(n17773), .D(n17772), .Y(n17781)
         );
  AOI22XL U21928 ( .A0(weight_1[294]), .A1(n17787), .B0(weight_1[270]), .B1(
        n17802), .Y(n17779) );
  AOI22XL U21929 ( .A0(weight_1[192]), .A1(n17884), .B0(weight_1[108]), .B1(
        n17792), .Y(n17778) );
  AOI22XL U21930 ( .A0(weight_1[120]), .A1(n17895), .B0(weight_1[12]), .B1(
        n17893), .Y(n17777) );
  AOI22XL U21931 ( .A0(weight_1[144]), .A1(n17868), .B0(weight_1[42]), .B1(
        n17789), .Y(n17776) );
  NAND4XL U21932 ( .A(n17779), .B(n17778), .C(n17777), .D(n17776), .Y(n17780)
         );
  NOR4XL U21933 ( .A(n17783), .B(n17782), .C(n17781), .D(n17780), .Y(n17784)
         );
  AOI32XL U21934 ( .A0(n17786), .A1(n17785), .A2(n17784), .B0(cursor[6]), .B1(
        n17785), .Y(n20647) );
  NAND2XL U21935 ( .A(n33554), .B(n20647), .Y(DP_OP_5168J1_124_9881_n57) );
  AOI22XL U21936 ( .A0(n21748), .A1(weight_1[301]), .B0(weight_1[295]), .B1(
        n17787), .Y(n17796) );
  AOI22XL U21937 ( .A0(n21999), .A1(weight_1[79]), .B0(weight_1[253]), .B1(
        n17788), .Y(n17795) );
  AOI22XL U21938 ( .A0(weight_1[175]), .A1(n17790), .B0(weight_1[43]), .B1(
        n17789), .Y(n17794) );
  AOI22XL U21939 ( .A0(weight_1[109]), .A1(n17792), .B0(weight_1[49]), .B1(
        n17791), .Y(n17793) );
  NAND4XL U21940 ( .A(n17796), .B(n17795), .C(n17794), .D(n17793), .Y(n17835)
         );
  AOI22XL U21941 ( .A0(weight_1[289]), .A1(n17798), .B0(weight_1[235]), .B1(
        n17797), .Y(n17808) );
  AOI22XL U21942 ( .A0(weight_1[379]), .A1(n17800), .B0(weight_1[67]), .B1(
        n17799), .Y(n17807) );
  AOI22XL U21943 ( .A0(weight_1[271]), .A1(n17802), .B0(weight_1[115]), .B1(
        n17801), .Y(n17806) );
  AOI22XL U21944 ( .A0(weight_1[205]), .A1(n17804), .B0(weight_1[37]), .B1(
        n17803), .Y(n17805) );
  NAND4XL U21945 ( .A(n17808), .B(n17807), .C(n17806), .D(n17805), .Y(n17834)
         );
  AOI22XL U21946 ( .A0(weight_1[367]), .A1(n17810), .B0(weight_1[361]), .B1(
        n17809), .Y(n17820) );
  AOI22XL U21947 ( .A0(weight_1[337]), .A1(n17812), .B0(weight_1[217]), .B1(
        n17811), .Y(n17819) );
  AOI22XL U21948 ( .A0(weight_1[325]), .A1(n17814), .B0(weight_1[187]), .B1(
        n17813), .Y(n17818) );
  AOI22XL U21949 ( .A0(weight_1[343]), .A1(n17816), .B0(weight_1[229]), .B1(
        n17815), .Y(n17817) );
  NAND4XL U21950 ( .A(n17820), .B(n17819), .C(n17818), .D(n17817), .Y(n17833)
         );
  AOI22XL U21951 ( .A0(n16744), .A1(weight_1[73]), .B0(weight_1[373]), .B1(
        n17821), .Y(n17831) );
  AOI22XL U21952 ( .A0(weight_1[331]), .A1(n17823), .B0(weight_1[139]), .B1(
        n17822), .Y(n17830) );
  AOI22XL U21953 ( .A0(weight_1[355]), .A1(n17825), .B0(weight_1[223]), .B1(
        n17824), .Y(n17829) );
  AOI22XL U21954 ( .A0(weight_1[349]), .A1(n17827), .B0(weight_1[283]), .B1(
        n17826), .Y(n17828) );
  NAND4XL U21955 ( .A(n17831), .B(n17830), .C(n17829), .D(n17828), .Y(n17832)
         );
  INVXL U21956 ( .A(weight_1[427]), .Y(n32421) );
  OAI22XL U21957 ( .A0(n32727), .A1(n17837), .B0(n32421), .B1(n17836), .Y(
        n17862) );
  INVXL U21958 ( .A(weight_1[421]), .Y(n32422) );
  INVXL U21959 ( .A(weight_1[385]), .Y(n32428) );
  OAI22XL U21960 ( .A0(n32422), .A1(n17839), .B0(n32428), .B1(n17838), .Y(
        n17861) );
  INVXL U21961 ( .A(weight_1[457]), .Y(n32419) );
  AOI22XL U21962 ( .A0(weight_1[481]), .A1(n17841), .B0(weight_1[403]), .B1(
        n17840), .Y(n17845) );
  AOI22XL U21963 ( .A0(weight_1[475]), .A1(n17843), .B0(weight_1[463]), .B1(
        n17842), .Y(n17844) );
  OAI211XL U21964 ( .A0(n32419), .A1(n17846), .B0(n17845), .C0(n17844), .Y(
        n17860) );
  AOI22XL U21965 ( .A0(weight_1[433]), .A1(n17848), .B0(weight_1[415]), .B1(
        n17847), .Y(n17858) );
  AOI22XL U21966 ( .A0(weight_1[469]), .A1(n17850), .B0(weight_1[439]), .B1(
        n17849), .Y(n17857) );
  AOI22XL U21967 ( .A0(weight_1[451]), .A1(n17852), .B0(weight_1[397]), .B1(
        n17851), .Y(n17856) );
  AOI22XL U21968 ( .A0(weight_1[409]), .A1(n17854), .B0(weight_1[391]), .B1(
        n17853), .Y(n17855) );
  NAND4XL U21969 ( .A(n17858), .B(n17857), .C(n17856), .D(n17855), .Y(n17859)
         );
  AOI22XL U21970 ( .A0(n26082), .A1(weight_1[313]), .B0(weight_1[151]), .B1(
        n17863), .Y(n17872) );
  AOI22XL U21971 ( .A0(n21766), .A1(weight_1[307]), .B0(weight_1[259]), .B1(
        n17864), .Y(n17871) );
  AOI22XL U21972 ( .A0(weight_1[181]), .A1(n17866), .B0(weight_1[61]), .B1(
        n17865), .Y(n17870) );
  AOI22XL U21973 ( .A0(weight_1[145]), .A1(n17868), .B0(weight_1[25]), .B1(
        n17867), .Y(n17869) );
  NAND4XL U21974 ( .A(n17872), .B(n17871), .C(n17870), .D(n17869), .Y(n17908)
         );
  AOI22XL U21975 ( .A0(weight_1[31]), .A1(n17874), .B0(weight_1[19]), .B1(
        n17873), .Y(n17882) );
  AOI22XL U21976 ( .A0(weight_1[169]), .A1(n16724), .B0(weight_1[133]), .B1(
        n17875), .Y(n17881) );
  AOI22XL U21977 ( .A0(weight_1[265]), .A1(n17877), .B0(weight_1[103]), .B1(
        n17876), .Y(n17880) );
  AOI22XL U21978 ( .A0(n26059), .A1(weight_1[319]), .B0(weight_1[211]), .B1(
        n17878), .Y(n17879) );
  NAND4XL U21979 ( .A(n17882), .B(n17881), .C(n17880), .D(n17879), .Y(n17907)
         );
  AOI22XL U21980 ( .A0(weight_1[193]), .A1(n17884), .B0(weight_1[55]), .B1(
        n17883), .Y(n17892) );
  AOI22XL U21981 ( .A0(weight_1[247]), .A1(n17886), .B0(weight_1[91]), .B1(
        n17885), .Y(n17891) );
  AOI22XL U21982 ( .A0(n21764), .A1(weight_1[7]), .B0(n21762), .B1(weight_1[1]), .Y(n17890) );
  AOI22XL U21983 ( .A0(weight_1[157]), .A1(n17888), .B0(weight_1[97]), .B1(
        n17887), .Y(n17889) );
  NAND4XL U21984 ( .A(n17892), .B(n17891), .C(n17890), .D(n17889), .Y(n17906)
         );
  AOI22XL U21985 ( .A0(weight_1[127]), .A1(n17894), .B0(weight_1[13]), .B1(
        n17893), .Y(n17904) );
  AOI22XL U21986 ( .A0(weight_1[241]), .A1(n17896), .B0(weight_1[121]), .B1(
        n17895), .Y(n17903) );
  AOI22XL U21987 ( .A0(weight_1[199]), .A1(n17898), .B0(weight_1[85]), .B1(
        n17897), .Y(n17902) );
  AOI22XL U21988 ( .A0(weight_1[277]), .A1(n17900), .B0(weight_1[163]), .B1(
        n17899), .Y(n17901) );
  NAND4XL U21989 ( .A(n17904), .B(n17903), .C(n17902), .D(n17901), .Y(n17905)
         );
  NAND2XL U21990 ( .A(n33554), .B(n20649), .Y(DP_OP_5168J1_124_9881_n56) );
  NAND2XL U21991 ( .A(n33068), .B(n20645), .Y(DP_OP_5168J1_124_9881_n76) );
  NAND2XL U21992 ( .A(n33554), .B(n20644), .Y(DP_OP_5168J1_124_9881_n55) );
  NAND2XL U21993 ( .A(n33554), .B(n17916), .Y(DP_OP_5168J1_124_9881_n54) );
  NAND2XL U21994 ( .A(n33068), .B(n17918), .Y(DP_OP_5168J1_124_9881_n58) );
  NAND2XL U21995 ( .A(n33554), .B(n17919), .Y(DP_OP_5168J1_124_9881_n53) );
  INVXL U21996 ( .A(affine_1[5]), .Y(DP_OP_5168J1_124_9881_n33) );
  AND2XL U21997 ( .A(n20649), .B(n20646), .Y(n17912) );
  AND2XL U21998 ( .A(n20649), .B(n17918), .Y(n17915) );
  AND2XL U21999 ( .A(n17916), .B(n20648), .Y(n17914) );
  ADDHXL U22000 ( .A(affine_1[3]), .B(n17912), .CO(n17913), .S(
        DP_OP_5168J1_124_9881_n45) );
  ADDFX1 U22001 ( .A(n17915), .B(n17914), .CI(n17913), .CO(
        DP_OP_5168J1_124_9881_n37), .S(DP_OP_5168J1_124_9881_n38) );
  AND2XL U22002 ( .A(n20645), .B(n17916), .Y(DP_OP_5168J1_124_9881_n78) );
  AND2XL U22003 ( .A(n17916), .B(n20646), .Y(DP_OP_5168J1_124_9881_n66) );
  AND2XL U22004 ( .A(n17919), .B(n20648), .Y(DP_OP_5168J1_124_9881_n71) );
  AND2XL U22005 ( .A(n17919), .B(n20646), .Y(DP_OP_5168J1_124_9881_n65) );
  AND2XL U22006 ( .A(n20647), .B(n17918), .Y(DP_OP_5168J1_124_9881_n63) );
  XOR2XL U22007 ( .A(affine_1[4]), .B(n17917), .Y(DP_OP_5168J1_124_9881_n40)
         );
  AND2XL U22008 ( .A(n17919), .B(n17918), .Y(n17921) );
  NAND2XL U22009 ( .A(n33068), .B(n20646), .Y(n17920) );
  AOI222XL U22010 ( .A0(counter[1]), .A1(affine_1[28]), .B0(n17988), .B1(
        affine_1[18]), .C0(n19228), .C1(affine_1[8]), .Y(n17922) );
  INVXL U22011 ( .A(weight_2[30]), .Y(n20413) );
  AOI22XL U22012 ( .A0(weight_2[48]), .A1(n17972), .B0(weight_2[12]), .B1(
        n18072), .Y(n17928) );
  INVXL U22013 ( .A(weight_2[24]), .Y(n20414) );
  INVXL U22014 ( .A(weight_2[18]), .Y(n20412) );
  OAI22XL U22015 ( .A0(n20414), .A1(n18118), .B0(n20412), .B1(n18117), .Y(
        n17926) );
  INVXL U22016 ( .A(weight_2[42]), .Y(n20417) );
  INVXL U22017 ( .A(weight_2[0]), .Y(n20393) );
  OAI22XL U22018 ( .A0(n20417), .A1(n18120), .B0(n20393), .B1(n17973), .Y(
        n17925) );
  INVXL U22019 ( .A(weight_2[36]), .Y(n20418) );
  INVXL U22020 ( .A(weight_2[6]), .Y(n20398) );
  OAI22XL U22021 ( .A0(n20418), .A1(n18127), .B0(n20398), .B1(n18043), .Y(
        n17924) );
  NOR3XL U22022 ( .A(n17926), .B(n17925), .C(n17924), .Y(n17927) );
  OAI211X1 U22023 ( .A0(n20413), .A1(n18109), .B0(n17928), .C0(n17927), .Y(
        n17929) );
  INVXL U22024 ( .A(weight_2[19]), .Y(n20408) );
  AOI22XL U22025 ( .A0(weight_2[49]), .A1(n17972), .B0(weight_2[13]), .B1(
        n18072), .Y(n17934) );
  INVXL U22026 ( .A(weight_2[31]), .Y(n20409) );
  INVXL U22027 ( .A(weight_2[25]), .Y(n20410) );
  OAI22XL U22028 ( .A0(n20409), .A1(n18109), .B0(n20410), .B1(n18118), .Y(
        n17932) );
  INVXL U22029 ( .A(weight_2[7]), .Y(n20403) );
  INVXL U22030 ( .A(weight_2[1]), .Y(n20402) );
  OAI22XL U22031 ( .A0(n20403), .A1(n18043), .B0(n20402), .B1(n17973), .Y(
        n17931) );
  INVXL U22032 ( .A(weight_2[43]), .Y(n20405) );
  INVXL U22033 ( .A(weight_2[37]), .Y(n20406) );
  OAI22XL U22034 ( .A0(n20405), .A1(n18120), .B0(n20406), .B1(n18127), .Y(
        n17930) );
  NOR3X1 U22035 ( .A(n17932), .B(n17931), .C(n17930), .Y(n17933) );
  OAI211XL U22036 ( .A0(n20408), .A1(n18117), .B0(n17934), .C0(n17933), .Y(
        n17935) );
  AOI222XL U22037 ( .A0(counter[1]), .A1(affine_1[29]), .B0(n17988), .B1(
        affine_1[19]), .C0(n19228), .C1(affine_1[9]), .Y(n17936) );
  MXI2XL U22038 ( .A(n19650), .B(n19647), .S0(n24570), .Y(n17937) );
  NAND2XL U22039 ( .A(n17929), .B(n17937), .Y(n17938) );
  OAI31XL U22040 ( .A0(n18151), .A1(n17929), .A2(n19650), .B0(n17938), .Y(
        n17939) );
  ADDHXL U22041 ( .A(affine_2[41]), .B(n17939), .CO(DP_OP_5169J1_125_4278_n40), 
        .S(DP_OP_5169J1_125_4278_n41) );
  AOI222XL U22042 ( .A0(counter[1]), .A1(affine_1[27]), .B0(n17988), .B1(
        affine_1[17]), .C0(n19228), .C1(affine_1[7]), .Y(n17940) );
  MXI2XL U22043 ( .A(n19647), .B(n19650), .S0(n18151), .Y(n17941) );
  OAI32XL U22044 ( .A0(n17929), .A1(n18149), .A2(n19650), .B0(n17941), .B1(
        n19651), .Y(n17942) );
  ADDHXL U22045 ( .A(affine_2[40]), .B(n17942), .CO(DP_OP_5169J1_125_4278_n45), 
        .S(DP_OP_5169J1_125_4278_n46) );
  AOI222XL U22046 ( .A0(counter[1]), .A1(affine_1[26]), .B0(n17988), .B1(
        affine_1[16]), .C0(n19228), .C1(affine_1[6]), .Y(n17943) );
  MXI2XL U22047 ( .A(n19647), .B(n19650), .S0(n18149), .Y(n17944) );
  OAI32XL U22048 ( .A0(n17929), .A1(n18147), .A2(n19650), .B0(n17944), .B1(
        n19651), .Y(n17945) );
  ADDHXL U22049 ( .A(affine_2[39]), .B(n17945), .CO(DP_OP_5169J1_125_4278_n50), 
        .S(DP_OP_5169J1_125_4278_n51) );
  AOI222XL U22050 ( .A0(counter[1]), .A1(affine_1[25]), .B0(n17988), .B1(
        affine_1[15]), .C0(n19228), .C1(affine_1[5]), .Y(n17946) );
  MXI2XL U22051 ( .A(n19647), .B(n19650), .S0(n18147), .Y(n17947) );
  OAI32XL U22052 ( .A0(n17929), .A1(n18145), .A2(n19650), .B0(n17947), .B1(
        n19651), .Y(n17948) );
  ADDHXL U22053 ( .A(affine_2[38]), .B(n17948), .CO(DP_OP_5169J1_125_4278_n55), 
        .S(DP_OP_5169J1_125_4278_n56) );
  AOI222XL U22054 ( .A0(counter[1]), .A1(affine_1[24]), .B0(n17988), .B1(
        affine_1[14]), .C0(n19228), .C1(affine_1[4]), .Y(n17949) );
  MXI2XL U22055 ( .A(n19647), .B(n19650), .S0(n18145), .Y(n17950) );
  OAI32XL U22056 ( .A0(n17929), .A1(n18141), .A2(n19650), .B0(n17950), .B1(
        n19651), .Y(n17951) );
  ADDHXL U22057 ( .A(affine_2[37]), .B(n17951), .CO(DP_OP_5169J1_125_4278_n60), 
        .S(DP_OP_5169J1_125_4278_n61) );
  AOI22XL U22058 ( .A0(weight_2[32]), .A1(n18115), .B0(weight_2[26]), .B1(
        n18108), .Y(n17956) );
  INVXL U22059 ( .A(n18127), .Y(n17971) );
  AOI22XL U22060 ( .A0(weight_2[50]), .A1(n17972), .B0(weight_2[38]), .B1(
        n17971), .Y(n17955) );
  INVXL U22061 ( .A(weight_2[44]), .Y(n20400) );
  INVXL U22062 ( .A(weight_2[8]), .Y(n20392) );
  OAI22XL U22063 ( .A0(n20400), .A1(n18120), .B0(n20392), .B1(n18043), .Y(
        n17953) );
  INVXL U22064 ( .A(weight_2[20]), .Y(n20395) );
  INVXL U22065 ( .A(weight_2[2]), .Y(n20391) );
  OAI22XL U22066 ( .A0(n20395), .A1(n18117), .B0(n20391), .B1(n17973), .Y(
        n17952) );
  AOI211XL U22067 ( .A0(weight_2[14]), .A1(n18072), .B0(n17953), .C0(n17952), 
        .Y(n17954) );
  NAND3X1 U22068 ( .A(n17956), .B(n17955), .C(n17954), .Y(n19636) );
  INVXL U22069 ( .A(weight_2[33]), .Y(n20385) );
  AOI22XL U22070 ( .A0(weight_2[51]), .A1(n17972), .B0(weight_2[15]), .B1(
        n18072), .Y(n17961) );
  INVXL U22071 ( .A(weight_2[27]), .Y(n20378) );
  INVXL U22072 ( .A(weight_2[21]), .Y(n20380) );
  OAI22XL U22073 ( .A0(n20378), .A1(n18118), .B0(n20380), .B1(n18117), .Y(
        n17959) );
  INVXL U22074 ( .A(weight_2[39]), .Y(n20388) );
  INVXL U22075 ( .A(weight_2[9]), .Y(n20383) );
  OAI22XL U22076 ( .A0(n20388), .A1(n18127), .B0(n20383), .B1(n18043), .Y(
        n17958) );
  INVXL U22077 ( .A(weight_2[45]), .Y(n20389) );
  INVXL U22078 ( .A(weight_2[3]), .Y(n20384) );
  OAI22XL U22079 ( .A0(n20389), .A1(n18120), .B0(n20384), .B1(n17973), .Y(
        n17957) );
  MXI2XL U22080 ( .A(n19638), .B(n17962), .S0(n18151), .Y(n17980) );
  INVXL U22081 ( .A(n19636), .Y(n17963) );
  MXI2XL U22082 ( .A(n19638), .B(n17962), .S0(n18149), .Y(n17981) );
  AOI22XL U22083 ( .A0(n19637), .A1(n17980), .B0(n18003), .B1(n17981), .Y(
        n18004) );
  NAND2BXL U22084 ( .AN(affine_2[42]), .B(n18004), .Y(
        DP_OP_5169J1_125_4278_n35) );
  INVXL U22085 ( .A(n18117), .Y(n17970) );
  AOI22XL U22086 ( .A0(weight_2[28]), .A1(n18108), .B0(weight_2[22]), .B1(
        n17970), .Y(n17968) );
  INVXL U22087 ( .A(weight_2[10]), .Y(n20386) );
  AOI2BB2XL U22088 ( .B0(weight_2[52]), .B1(n17972), .A0N(n20386), .A1N(n18043), .Y(n17967) );
  INVXL U22089 ( .A(weight_2[46]), .Y(n20370) );
  INVXL U22090 ( .A(weight_2[40]), .Y(n20371) );
  OAI22XL U22091 ( .A0(n20370), .A1(n18120), .B0(n20371), .B1(n18127), .Y(
        n17965) );
  INVXL U22092 ( .A(weight_2[16]), .Y(n20376) );
  INVXL U22093 ( .A(weight_2[4]), .Y(n20387) );
  OAI22XL U22094 ( .A0(n20376), .A1(n18116), .B0(n20387), .B1(n17973), .Y(
        n17964) );
  AOI211XL U22095 ( .A0(weight_2[34]), .A1(n18115), .B0(n17965), .C0(n17964), 
        .Y(n17966) );
  MXI2X1 U22096 ( .A(n19638), .B(n17962), .S0(n17983), .Y(n24545) );
  INVX2 U22097 ( .A(n24545), .Y(n28211) );
  AOI22XL U22098 ( .A0(weight_2[23]), .A1(n17970), .B0(weight_2[17]), .B1(
        n18072), .Y(n17978) );
  AOI22XL U22099 ( .A0(weight_2[53]), .A1(n17972), .B0(weight_2[41]), .B1(
        n17971), .Y(n17977) );
  INVXL U22100 ( .A(weight_2[47]), .Y(n20377) );
  INVXL U22101 ( .A(weight_2[11]), .Y(n20369) );
  OAI22XL U22102 ( .A0(n20377), .A1(n18120), .B0(n20369), .B1(n18043), .Y(
        n17975) );
  INVXL U22103 ( .A(weight_2[29]), .Y(n20365) );
  INVXL U22104 ( .A(weight_2[5]), .Y(n20367) );
  OAI22XL U22105 ( .A0(n20365), .A1(n18118), .B0(n20367), .B1(n17973), .Y(
        n17974) );
  AOI211XL U22106 ( .A0(weight_2[35]), .A1(n18115), .B0(n17975), .C0(n17974), 
        .Y(n17976) );
  INVX1 U22107 ( .A(n24543), .Y(n24544) );
  AOI221XL U22108 ( .A0(n24545), .A1(n19698), .B0(n28211), .B1(n17983), .C0(
        n24544), .Y(DP_OP_5169J1_125_4278_n76) );
  MXI2XL U22109 ( .A(n19638), .B(n17962), .S0(n24570), .Y(n18002) );
  NAND2XL U22110 ( .A(n18002), .B(n19637), .Y(n17979) );
  OAI2BB1XL U22111 ( .A0N(n17980), .A1N(n18003), .B0(n17979), .Y(
        DP_OP_5169J1_125_4278_n91) );
  MXI2XL U22112 ( .A(n17962), .B(n19638), .S0(n18147), .Y(n17998) );
  OAI2BB2XL U22113 ( .B0(n19640), .B1(n17998), .A0N(n19637), .A1N(n17981), .Y(
        DP_OP_5169J1_125_4278_n93) );
  AOI222XL U22114 ( .A0(counter[1]), .A1(affine_1[21]), .B0(n17988), .B1(
        affine_1[11]), .C0(n19228), .C1(affine_1[1]), .Y(n17982) );
  INVXL U22115 ( .A(n17982), .Y(n19666) );
  MXI2XL U22116 ( .A(n24543), .B(n24544), .S0(n19666), .Y(n17987) );
  INVXL U22117 ( .A(n17983), .Y(n17984) );
  AOI22XL U22118 ( .A0(n19698), .A1(n24544), .B0(n24543), .B1(n19652), .Y(
        n17985) );
  OAI22XL U22119 ( .A0(n28211), .A1(n17987), .B0(n28210), .B1(n17985), .Y(
        DP_OP_5169J1_125_4278_n88) );
  INVX1 U22120 ( .A(n19637), .Y(n19643) );
  AOI222XL U22121 ( .A0(counter[1]), .A1(affine_1[22]), .B0(n17988), .B1(
        affine_1[12]), .C0(n19228), .C1(affine_1[2]), .Y(n17986) );
  INVXL U22122 ( .A(n17986), .Y(n19694) );
  MXI2XL U22123 ( .A(n17962), .B(n19638), .S0(n19694), .Y(n17990) );
  MXI2XL U22124 ( .A(n17962), .B(n19638), .S0(n19666), .Y(n19641) );
  OAI22XL U22125 ( .A0(n19643), .A1(n17990), .B0(n19640), .B1(n19641), .Y(
        DP_OP_5169J1_125_4278_n98) );
  MXI2XL U22126 ( .A(n24543), .B(n24544), .S0(n19694), .Y(n17992) );
  OAI22XL U22127 ( .A0(n28211), .A1(n17992), .B0(n28210), .B1(n17987), .Y(
        DP_OP_5169J1_125_4278_n87) );
  AOI222XL U22128 ( .A0(counter[1]), .A1(affine_1[23]), .B0(n17988), .B1(
        affine_1[13]), .C0(n19228), .C1(affine_1[3]), .Y(n17989) );
  MXI2XL U22129 ( .A(n17962), .B(n19638), .S0(n19689), .Y(n17993) );
  OAI22XL U22130 ( .A0(n19643), .A1(n17993), .B0(n19640), .B1(n17990), .Y(
        DP_OP_5169J1_125_4278_n97) );
  MXI2XL U22131 ( .A(n19647), .B(n19650), .S0(n18141), .Y(n17991) );
  OAI32XL U22132 ( .A0(n17929), .A1(n19689), .A2(n19650), .B0(n17991), .B1(
        n19651), .Y(DP_OP_5169J1_125_4278_n107) );
  MXI2XL U22133 ( .A(n24543), .B(n24544), .S0(n19689), .Y(n17994) );
  OAI22XL U22134 ( .A0(n28211), .A1(n17994), .B0(n28210), .B1(n17992), .Y(
        DP_OP_5169J1_125_4278_n86) );
  MXI2XL U22135 ( .A(n17962), .B(n19638), .S0(n18141), .Y(n17995) );
  OAI22XL U22136 ( .A0(n19643), .A1(n17995), .B0(n19640), .B1(n17993), .Y(
        DP_OP_5169J1_125_4278_n96) );
  MXI2XL U22137 ( .A(n24543), .B(n24544), .S0(n18141), .Y(n17996) );
  OAI22XL U22138 ( .A0(n28211), .A1(n17996), .B0(n28210), .B1(n17994), .Y(
        DP_OP_5169J1_125_4278_n85) );
  MXI2XL U22139 ( .A(n17962), .B(n19638), .S0(n18145), .Y(n17997) );
  OAI22XL U22140 ( .A0(n19643), .A1(n17997), .B0(n19640), .B1(n17995), .Y(
        DP_OP_5169J1_125_4278_n95) );
  MXI2XL U22141 ( .A(n24543), .B(n24544), .S0(n18145), .Y(n17999) );
  OAI22XL U22142 ( .A0(n28211), .A1(n17999), .B0(n28210), .B1(n17996), .Y(
        DP_OP_5169J1_125_4278_n84) );
  OAI22XL U22143 ( .A0(n19643), .A1(n17998), .B0(n19640), .B1(n17997), .Y(
        DP_OP_5169J1_125_4278_n94) );
  MXI2XL U22144 ( .A(n24543), .B(n24544), .S0(n18147), .Y(n18000) );
  OAI22XL U22145 ( .A0(n28211), .A1(n18000), .B0(n28210), .B1(n17999), .Y(
        DP_OP_5169J1_125_4278_n83) );
  MXI2XL U22146 ( .A(n24543), .B(n24544), .S0(n18149), .Y(n18001) );
  OAI22XL U22147 ( .A0(n28211), .A1(n18001), .B0(n28210), .B1(n18000), .Y(
        DP_OP_5169J1_125_4278_n82) );
  MXI2XL U22148 ( .A(n24543), .B(n24544), .S0(n18151), .Y(n24546) );
  OAI22XL U22149 ( .A0(n28211), .A1(n24546), .B0(n28210), .B1(n18001), .Y(
        DP_OP_5169J1_125_4278_n81) );
  AOI32XL U22150 ( .A0(n17929), .A1(n24570), .A2(n19650), .B0(n19647), .B1(
        n17936), .Y(DP_OP_5169J1_125_4278_n101) );
  OAI21XL U22151 ( .A0(n19637), .A1(n18003), .B0(n18002), .Y(
        DP_OP_5169J1_125_4278_n90) );
  INVXL U22152 ( .A(affine_2[43]), .Y(DP_OP_5169J1_125_4278_n31) );
  XOR2XL U22153 ( .A(affine_2[42]), .B(n18004), .Y(DP_OP_5169J1_125_4278_n36)
         );
  OAI22XL U22154 ( .A0(n20418), .A1(n18120), .B0(n20413), .B1(n18127), .Y(
        n18008) );
  NAND2X2 U22155 ( .A(n19097), .B(n19221), .Y(n18121) );
  OAI22XL U22156 ( .A0(n20417), .A1(n18121), .B0(n20393), .B1(n18043), .Y(
        n18007) );
  INVXL U22157 ( .A(weight_2[12]), .Y(n20411) );
  OAI22XL U22158 ( .A0(n20411), .A1(n18117), .B0(n20398), .B1(n18116), .Y(
        n18006) );
  OAI22XL U22159 ( .A0(n20414), .A1(n18109), .B0(n20412), .B1(n18118), .Y(
        n18005) );
  NOR4XL U22160 ( .A(n18008), .B(n18007), .C(n18006), .D(n18005), .Y(n18009)
         );
  OAI22XL U22161 ( .A0(n20405), .A1(n18121), .B0(n20409), .B1(n18127), .Y(
        n18014) );
  OAI22XL U22162 ( .A0(n20406), .A1(n18120), .B0(n20402), .B1(n18043), .Y(
        n18013) );
  OAI22XL U22163 ( .A0(n20408), .A1(n18118), .B0(n20403), .B1(n18116), .Y(
        n18012) );
  INVXL U22164 ( .A(weight_2[13]), .Y(n20407) );
  OAI22XL U22165 ( .A0(n20410), .A1(n18109), .B0(n20407), .B1(n18117), .Y(
        n18011) );
  MXI2XL U22166 ( .A(n19629), .B(n19626), .S0(n24570), .Y(n18016) );
  NAND2XL U22167 ( .A(n18010), .B(n18016), .Y(n18017) );
  OAI31XL U22168 ( .A0(n18151), .A1(n18010), .A2(n19629), .B0(n18017), .Y(
        n18018) );
  ADDHXL U22169 ( .A(affine_2[25]), .B(n18018), .CO(DP_OP_5170J1_126_4278_n40), 
        .S(DP_OP_5170J1_126_4278_n41) );
  MXI2XL U22170 ( .A(n19626), .B(n19629), .S0(n18151), .Y(n18019) );
  OAI32XL U22171 ( .A0(n18010), .A1(n18149), .A2(n19629), .B0(n18019), .B1(
        n19630), .Y(n18020) );
  ADDHXL U22172 ( .A(affine_2[24]), .B(n18020), .CO(DP_OP_5170J1_126_4278_n45), 
        .S(DP_OP_5170J1_126_4278_n46) );
  MXI2XL U22173 ( .A(n19626), .B(n19629), .S0(n18149), .Y(n18021) );
  OAI32XL U22174 ( .A0(n18010), .A1(n18147), .A2(n19629), .B0(n18021), .B1(
        n19630), .Y(n18022) );
  ADDHXL U22175 ( .A(affine_2[23]), .B(n18022), .CO(DP_OP_5170J1_126_4278_n50), 
        .S(DP_OP_5170J1_126_4278_n51) );
  MXI2XL U22176 ( .A(n19626), .B(n19629), .S0(n18147), .Y(n18023) );
  OAI32XL U22177 ( .A0(n18010), .A1(n18145), .A2(n19629), .B0(n18023), .B1(
        n19630), .Y(n18024) );
  ADDHXL U22178 ( .A(affine_2[22]), .B(n18024), .CO(DP_OP_5170J1_126_4278_n55), 
        .S(DP_OP_5170J1_126_4278_n56) );
  MXI2XL U22179 ( .A(n19626), .B(n19629), .S0(n18145), .Y(n18025) );
  OAI32XL U22180 ( .A0(n18010), .A1(n18141), .A2(n19629), .B0(n18025), .B1(
        n19630), .Y(n18026) );
  ADDHXL U22181 ( .A(affine_2[21]), .B(n18026), .CO(DP_OP_5170J1_126_4278_n60), 
        .S(DP_OP_5170J1_126_4278_n61) );
  INVXL U22182 ( .A(weight_2[32]), .Y(n20396) );
  OAI22XL U22183 ( .A0(n20396), .A1(n18127), .B0(n20391), .B1(n18043), .Y(
        n18030) );
  INVXL U22184 ( .A(weight_2[38]), .Y(n20399) );
  OAI22XL U22185 ( .A0(n20400), .A1(n18121), .B0(n20399), .B1(n18120), .Y(
        n18029) );
  INVXL U22186 ( .A(weight_2[14]), .Y(n20394) );
  OAI22XL U22187 ( .A0(n20394), .A1(n18117), .B0(n20392), .B1(n18116), .Y(
        n18028) );
  INVXL U22188 ( .A(weight_2[26]), .Y(n20397) );
  OAI22XL U22189 ( .A0(n20397), .A1(n18109), .B0(n20395), .B1(n18118), .Y(
        n18027) );
  NOR4XL U22190 ( .A(n18030), .B(n18029), .C(n18028), .D(n18027), .Y(n18031)
         );
  OAI22XL U22191 ( .A0(n20389), .A1(n18121), .B0(n20385), .B1(n18127), .Y(
        n18035) );
  OAI22XL U22192 ( .A0(n20388), .A1(n18120), .B0(n20384), .B1(n18043), .Y(
        n18034) );
  OAI22XL U22193 ( .A0(n20380), .A1(n18118), .B0(n20383), .B1(n18116), .Y(
        n18033) );
  INVXL U22194 ( .A(weight_2[15]), .Y(n20381) );
  OAI22XL U22195 ( .A0(n20378), .A1(n18109), .B0(n20381), .B1(n18117), .Y(
        n18032) );
  INVX1 U22196 ( .A(n19614), .Y(n19613) );
  MXI2XL U22197 ( .A(n19613), .B(n19614), .S0(n18151), .Y(n18051) );
  INVXL U22198 ( .A(n19611), .Y(n18037) );
  MXI2XL U22199 ( .A(n19613), .B(n19614), .S0(n18149), .Y(n18052) );
  AOI22XL U22200 ( .A0(n19612), .A1(n18051), .B0(n18070), .B1(n18052), .Y(
        n18071) );
  NAND2BXL U22201 ( .AN(affine_2[26]), .B(n18071), .Y(
        DP_OP_5170J1_126_4278_n35) );
  OAI22XL U22202 ( .A0(n20370), .A1(n18121), .B0(n20387), .B1(n18043), .Y(
        n18041) );
  INVXL U22203 ( .A(weight_2[34]), .Y(n20372) );
  OAI22XL U22204 ( .A0(n20371), .A1(n18120), .B0(n20372), .B1(n18127), .Y(
        n18040) );
  INVXL U22205 ( .A(weight_2[22]), .Y(n20374) );
  OAI22XL U22206 ( .A0(n20374), .A1(n18118), .B0(n20386), .B1(n18116), .Y(
        n18039) );
  INVXL U22207 ( .A(weight_2[28]), .Y(n20373) );
  OAI22XL U22208 ( .A0(n20373), .A1(n18109), .B0(n20376), .B1(n18117), .Y(
        n18038) );
  NOR4XL U22209 ( .A(n18041), .B(n18040), .C(n18039), .D(n18038), .Y(n18042)
         );
  OAI22XL U22210 ( .A0(n20377), .A1(n18121), .B0(n20367), .B1(n18043), .Y(
        n18047) );
  INVXL U22211 ( .A(weight_2[41]), .Y(n20375) );
  INVXL U22212 ( .A(weight_2[35]), .Y(n20364) );
  OAI22XL U22213 ( .A0(n20375), .A1(n18120), .B0(n20364), .B1(n18127), .Y(
        n18046) );
  INVXL U22214 ( .A(weight_2[23]), .Y(n20366) );
  OAI22XL U22215 ( .A0(n20365), .A1(n18109), .B0(n20366), .B1(n18118), .Y(
        n18045) );
  INVXL U22216 ( .A(weight_2[17]), .Y(n20368) );
  OAI22XL U22217 ( .A0(n20368), .A1(n18117), .B0(n20369), .B1(n18116), .Y(
        n18044) );
  NOR4XL U22218 ( .A(n18047), .B(n18046), .C(n18045), .D(n18044), .Y(n18048)
         );
  AOI221XL U22219 ( .A0(n24562), .A1(n19698), .B0(n28398), .B1(n18053), .C0(
        n24561), .Y(DP_OP_5170J1_126_4278_n76) );
  MXI2XL U22220 ( .A(n19613), .B(n19614), .S0(n24570), .Y(n18069) );
  NAND2XL U22221 ( .A(n18069), .B(n19612), .Y(n18050) );
  OAI2BB1XL U22222 ( .A0N(n18051), .A1N(n18070), .B0(n18050), .Y(
        DP_OP_5170J1_126_4278_n91) );
  MXI2XL U22223 ( .A(n19614), .B(n19613), .S0(n18147), .Y(n18064) );
  OAI2BB2XL U22224 ( .B0(n19616), .B1(n18064), .A0N(n19612), .A1N(n18052), .Y(
        DP_OP_5170J1_126_4278_n93) );
  MXI2XL U22225 ( .A(n19614), .B(n19613), .S0(n19694), .Y(n18056) );
  MXI2XL U22226 ( .A(n19614), .B(n19613), .S0(n19666), .Y(n19617) );
  OAI22XL U22227 ( .A0(n19622), .A1(n18056), .B0(n19616), .B1(n19617), .Y(
        DP_OP_5170J1_126_4278_n98) );
  INVXL U22228 ( .A(n18053), .Y(n18054) );
  AOI22XL U22229 ( .A0(n19698), .A1(n24561), .B0(n24560), .B1(n17969), .Y(
        n18055) );
  OAI22XL U22230 ( .A0(n28398), .A1(n18057), .B0(n28397), .B1(n18055), .Y(
        DP_OP_5170J1_126_4278_n88) );
  MXI2XL U22231 ( .A(n19614), .B(n19613), .S0(n19689), .Y(n18060) );
  OAI22XL U22232 ( .A0(n19622), .A1(n18060), .B0(n19616), .B1(n18056), .Y(
        DP_OP_5170J1_126_4278_n97) );
  OAI22XL U22233 ( .A0(n28398), .A1(n18059), .B0(n28397), .B1(n18057), .Y(
        DP_OP_5170J1_126_4278_n87) );
  MXI2XL U22234 ( .A(n19626), .B(n19629), .S0(n18141), .Y(n18058) );
  OAI32XL U22235 ( .A0(n18010), .A1(n19689), .A2(n19629), .B0(n18058), .B1(
        n19630), .Y(DP_OP_5170J1_126_4278_n107) );
  MXI2XL U22236 ( .A(n24560), .B(n24561), .S0(n19689), .Y(n18062) );
  OAI22XL U22237 ( .A0(n28398), .A1(n18062), .B0(n28397), .B1(n18059), .Y(
        DP_OP_5170J1_126_4278_n86) );
  MXI2XL U22238 ( .A(n19614), .B(n19613), .S0(n18141), .Y(n18061) );
  OAI22XL U22239 ( .A0(n19622), .A1(n18061), .B0(n19616), .B1(n18060), .Y(
        DP_OP_5170J1_126_4278_n96) );
  MXI2XL U22240 ( .A(n19614), .B(n19613), .S0(n18145), .Y(n18063) );
  OAI22XL U22241 ( .A0(n19622), .A1(n18063), .B0(n19616), .B1(n18061), .Y(
        DP_OP_5170J1_126_4278_n95) );
  MXI2XL U22242 ( .A(n24560), .B(n24561), .S0(n18141), .Y(n18065) );
  OAI22XL U22243 ( .A0(n28398), .A1(n18065), .B0(n28397), .B1(n18062), .Y(
        DP_OP_5170J1_126_4278_n85) );
  OAI22XL U22244 ( .A0(n19622), .A1(n18064), .B0(n19616), .B1(n18063), .Y(
        DP_OP_5170J1_126_4278_n94) );
  MXI2XL U22245 ( .A(n24560), .B(n24561), .S0(n18145), .Y(n18066) );
  OAI22XL U22246 ( .A0(n28398), .A1(n18066), .B0(n28397), .B1(n18065), .Y(
        DP_OP_5170J1_126_4278_n84) );
  MXI2XL U22247 ( .A(n24560), .B(n24561), .S0(n18147), .Y(n18067) );
  OAI22XL U22248 ( .A0(n28398), .A1(n18067), .B0(n28397), .B1(n18066), .Y(
        DP_OP_5170J1_126_4278_n83) );
  MXI2XL U22249 ( .A(n24560), .B(n24561), .S0(n18149), .Y(n18068) );
  OAI22XL U22250 ( .A0(n28398), .A1(n18068), .B0(n28397), .B1(n18067), .Y(
        DP_OP_5170J1_126_4278_n82) );
  MXI2XL U22251 ( .A(n24560), .B(n24561), .S0(n18151), .Y(n24563) );
  OAI22XL U22252 ( .A0(n28398), .A1(n24563), .B0(n28397), .B1(n18068), .Y(
        DP_OP_5170J1_126_4278_n81) );
  AOI32XL U22253 ( .A0(n18010), .A1(n24570), .A2(n19629), .B0(n19626), .B1(
        n17936), .Y(DP_OP_5170J1_126_4278_n101) );
  OAI21XL U22254 ( .A0(n19612), .A1(n18070), .B0(n18069), .Y(
        DP_OP_5170J1_126_4278_n90) );
  INVXL U22255 ( .A(affine_2[27]), .Y(DP_OP_5170J1_126_4278_n31) );
  XOR2XL U22256 ( .A(affine_2[26]), .B(n18071), .Y(DP_OP_5170J1_126_4278_n36)
         );
  AOI22XL U22257 ( .A0(N18014), .A1(weight_2[48]), .B0(weight_2[0]), .B1(
        n18072), .Y(n18077) );
  OAI22XL U22258 ( .A0(n20412), .A1(n18109), .B0(n20398), .B1(n18117), .Y(
        n18075) );
  OAI22XL U22259 ( .A0(n20418), .A1(n18121), .B0(n20411), .B1(n18118), .Y(
        n18074) );
  OAI22XL U22260 ( .A0(n20417), .A1(n18119), .B0(n20413), .B1(n18120), .Y(
        n18073) );
  NOR3XL U22261 ( .A(n18075), .B(n18074), .C(n18073), .Y(n18076) );
  OAI211X1 U22262 ( .A0(n20414), .A1(n18127), .B0(n18077), .C0(n18076), .Y(
        n18078) );
  AOI22XL U22263 ( .A0(N18014), .A1(weight_2[49]), .B0(weight_2[13]), .B1(
        n18108), .Y(n18083) );
  OAI22XL U22264 ( .A0(n20408), .A1(n18109), .B0(n20402), .B1(n18116), .Y(
        n18081) );
  OAI22XL U22265 ( .A0(n20410), .A1(n18127), .B0(n20403), .B1(n18117), .Y(
        n18080) );
  OAI22XL U22266 ( .A0(n20406), .A1(n18121), .B0(n20409), .B1(n18120), .Y(
        n18079) );
  NOR3X1 U22267 ( .A(n18081), .B(n18080), .C(n18079), .Y(n18082) );
  INVX3 U22268 ( .A(n18084), .Y(n19693) );
  MXI2XL U22269 ( .A(n19693), .B(n18084), .S0(n24570), .Y(n18085) );
  NAND2XL U22270 ( .A(n18078), .B(n18085), .Y(n18086) );
  OAI31XL U22271 ( .A0(n18151), .A1(n18078), .A2(n19693), .B0(n18086), .Y(
        n18087) );
  ADDHXL U22272 ( .A(affine_2[9]), .B(n18087), .CO(DP_OP_5171J1_127_4278_n40), 
        .S(DP_OP_5171J1_127_4278_n41) );
  MXI2XL U22273 ( .A(n18084), .B(n19693), .S0(n18151), .Y(n18088) );
  OAI32XL U22274 ( .A0(n18078), .A1(n18149), .A2(n19693), .B0(n18088), .B1(
        n19691), .Y(n18089) );
  ADDHXL U22275 ( .A(affine_2[8]), .B(n18089), .CO(DP_OP_5171J1_127_4278_n45), 
        .S(DP_OP_5171J1_127_4278_n46) );
  MXI2XL U22276 ( .A(n18084), .B(n19693), .S0(n18149), .Y(n18090) );
  OAI32XL U22277 ( .A0(n18078), .A1(n18147), .A2(n19693), .B0(n18090), .B1(
        n19691), .Y(n18091) );
  ADDHXL U22278 ( .A(affine_2[7]), .B(n18091), .CO(DP_OP_5171J1_127_4278_n50), 
        .S(DP_OP_5171J1_127_4278_n51) );
  MXI2XL U22279 ( .A(n18084), .B(n19693), .S0(n18147), .Y(n18092) );
  OAI32XL U22280 ( .A0(n18078), .A1(n18145), .A2(n19693), .B0(n18092), .B1(
        n19691), .Y(n18093) );
  ADDHXL U22281 ( .A(affine_2[6]), .B(n18093), .CO(DP_OP_5171J1_127_4278_n55), 
        .S(DP_OP_5171J1_127_4278_n56) );
  MXI2XL U22282 ( .A(n18084), .B(n19693), .S0(n18145), .Y(n18094) );
  OAI32XL U22283 ( .A0(n18078), .A1(n18141), .A2(n19693), .B0(n18094), .B1(
        n19691), .Y(n18095) );
  ADDHXL U22284 ( .A(affine_2[5]), .B(n18095), .CO(DP_OP_5171J1_127_4278_n60), 
        .S(DP_OP_5171J1_127_4278_n61) );
  AOI22XL U22285 ( .A0(N18014), .A1(weight_2[50]), .B0(weight_2[20]), .B1(
        n18115), .Y(n18100) );
  OAI22XL U22286 ( .A0(n20392), .A1(n18117), .B0(n20391), .B1(n18116), .Y(
        n18098) );
  OAI22XL U22287 ( .A0(n20400), .A1(n18119), .B0(n20394), .B1(n18118), .Y(
        n18097) );
  OAI22XL U22288 ( .A0(n20399), .A1(n18121), .B0(n20396), .B1(n18120), .Y(
        n18096) );
  MXI2X1 U22289 ( .A(n19693), .B(n18084), .S0(n19695), .Y(n19696) );
  AOI22XL U22290 ( .A0(N18014), .A1(weight_2[51]), .B0(weight_2[15]), .B1(
        n18108), .Y(n18105) );
  OAI22XL U22291 ( .A0(n20383), .A1(n18117), .B0(n20384), .B1(n18116), .Y(
        n18103) );
  OAI22XL U22292 ( .A0(n20385), .A1(n18120), .B0(n20380), .B1(n18109), .Y(
        n18102) );
  OAI22XL U22293 ( .A0(n20388), .A1(n18121), .B0(n20378), .B1(n18127), .Y(
        n18101) );
  MXI2XL U22294 ( .A(n19697), .B(n18106), .S0(n18151), .Y(n18130) );
  INVXL U22295 ( .A(n19695), .Y(n18107) );
  MXI2XL U22296 ( .A(n19697), .B(n18106), .S0(n18149), .Y(n18131) );
  AOI22XL U22297 ( .A0(n19696), .A1(n18130), .B0(n18154), .B1(n18131), .Y(
        n18155) );
  NAND2BXL U22298 ( .AN(affine_2[10]), .B(n18155), .Y(
        DP_OP_5171J1_127_4278_n35) );
  AOI22XL U22299 ( .A0(N18014), .A1(weight_2[52]), .B0(weight_2[16]), .B1(
        n18108), .Y(n18114) );
  OAI22XL U22300 ( .A0(n20374), .A1(n18109), .B0(n20387), .B1(n18116), .Y(
        n18112) );
  OAI22XL U22301 ( .A0(n20370), .A1(n18119), .B0(n20386), .B1(n18117), .Y(
        n18111) );
  OAI22XL U22302 ( .A0(n20372), .A1(n18120), .B0(n20373), .B1(n18127), .Y(
        n18110) );
  NOR3XL U22303 ( .A(n18112), .B(n18111), .C(n18110), .Y(n18113) );
  MXI2X1 U22304 ( .A(n19697), .B(n18106), .S0(n18132), .Y(n24572) );
  AOI22XL U22305 ( .A0(N18014), .A1(weight_2[53]), .B0(weight_2[23]), .B1(
        n18115), .Y(n18126) );
  OAI22XL U22306 ( .A0(n20369), .A1(n18117), .B0(n20367), .B1(n18116), .Y(
        n18124) );
  OAI22XL U22307 ( .A0(n20377), .A1(n18119), .B0(n20368), .B1(n18118), .Y(
        n18123) );
  OAI22XL U22308 ( .A0(n20375), .A1(n18121), .B0(n20364), .B1(n18120), .Y(
        n18122) );
  NOR3XL U22309 ( .A(n18124), .B(n18123), .C(n18122), .Y(n18125) );
  AOI221XL U22310 ( .A0(n24572), .A1(n19698), .B0(n28611), .B1(n18132), .C0(
        n24571), .Y(DP_OP_5171J1_127_4278_n76) );
  MXI2XL U22311 ( .A(n19697), .B(n18106), .S0(n24570), .Y(n18153) );
  NAND2XL U22312 ( .A(n18153), .B(n19696), .Y(n18129) );
  OAI2BB1XL U22313 ( .A0N(n18130), .A1N(n18154), .B0(n18129), .Y(
        DP_OP_5171J1_127_4278_n91) );
  INVX2 U22314 ( .A(n18154), .Y(n19701) );
  MXI2XL U22315 ( .A(n18106), .B(n19697), .S0(n18147), .Y(n18144) );
  OAI2BB2XL U22316 ( .B0(n19701), .B1(n18144), .A0N(n19696), .A1N(n18131), .Y(
        DP_OP_5171J1_127_4278_n93) );
  INVX1 U22317 ( .A(n19696), .Y(n19703) );
  MXI2XL U22318 ( .A(n18106), .B(n19697), .S0(n19694), .Y(n18135) );
  MXI2XL U22319 ( .A(n18106), .B(n19697), .S0(n19666), .Y(n19702) );
  OAI22XL U22320 ( .A0(n19703), .A1(n18135), .B0(n19701), .B1(n19702), .Y(
        DP_OP_5171J1_127_4278_n98) );
  MXI2XL U22321 ( .A(n18128), .B(n24571), .S0(n19666), .Y(n18136) );
  INVXL U22322 ( .A(n18132), .Y(n18133) );
  AOI22XL U22323 ( .A0(n19698), .A1(n24571), .B0(n18128), .B1(n17969), .Y(
        n18134) );
  OAI22XL U22324 ( .A0(n28611), .A1(n18136), .B0(n28610), .B1(n18134), .Y(
        DP_OP_5171J1_127_4278_n88) );
  MXI2XL U22325 ( .A(n18106), .B(n19697), .S0(n19689), .Y(n18139) );
  OAI22XL U22326 ( .A0(n19703), .A1(n18139), .B0(n19701), .B1(n18135), .Y(
        DP_OP_5171J1_127_4278_n97) );
  MXI2XL U22327 ( .A(n18128), .B(n24571), .S0(n19694), .Y(n18138) );
  OAI22XL U22328 ( .A0(n28611), .A1(n18138), .B0(n28610), .B1(n18136), .Y(
        DP_OP_5171J1_127_4278_n87) );
  MXI2XL U22329 ( .A(n18084), .B(n19693), .S0(n18141), .Y(n18137) );
  OAI32XL U22330 ( .A0(n18078), .A1(n19689), .A2(n19693), .B0(n18137), .B1(
        n19691), .Y(DP_OP_5171J1_127_4278_n107) );
  MXI2XL U22331 ( .A(n18128), .B(n24571), .S0(n19689), .Y(n18142) );
  OAI22XL U22332 ( .A0(n28611), .A1(n18142), .B0(n28610), .B1(n18138), .Y(
        DP_OP_5171J1_127_4278_n86) );
  MXI2XL U22333 ( .A(n18106), .B(n19697), .S0(n18141), .Y(n18140) );
  OAI22XL U22334 ( .A0(n19703), .A1(n18140), .B0(n19701), .B1(n18139), .Y(
        DP_OP_5171J1_127_4278_n96) );
  MXI2XL U22335 ( .A(n18106), .B(n19697), .S0(n18145), .Y(n18143) );
  OAI22XL U22336 ( .A0(n19703), .A1(n18143), .B0(n19701), .B1(n18140), .Y(
        DP_OP_5171J1_127_4278_n95) );
  MXI2XL U22337 ( .A(n18128), .B(n24571), .S0(n18141), .Y(n18146) );
  OAI22XL U22338 ( .A0(n28611), .A1(n18146), .B0(n28610), .B1(n18142), .Y(
        DP_OP_5171J1_127_4278_n85) );
  OAI22XL U22339 ( .A0(n19703), .A1(n18144), .B0(n19701), .B1(n18143), .Y(
        DP_OP_5171J1_127_4278_n94) );
  MXI2XL U22340 ( .A(n18128), .B(n24571), .S0(n18145), .Y(n18148) );
  OAI22XL U22341 ( .A0(n28611), .A1(n18148), .B0(n28610), .B1(n18146), .Y(
        DP_OP_5171J1_127_4278_n84) );
  MXI2XL U22342 ( .A(n18128), .B(n24571), .S0(n18147), .Y(n18150) );
  OAI22XL U22343 ( .A0(n28611), .A1(n18150), .B0(n28610), .B1(n18148), .Y(
        DP_OP_5171J1_127_4278_n83) );
  MXI2XL U22344 ( .A(n18128), .B(n24571), .S0(n18149), .Y(n18152) );
  OAI22XL U22345 ( .A0(n28611), .A1(n18152), .B0(n28610), .B1(n18150), .Y(
        DP_OP_5171J1_127_4278_n82) );
  MXI2XL U22346 ( .A(n18128), .B(n24571), .S0(n18151), .Y(n24573) );
  OAI22XL U22347 ( .A0(n28611), .A1(n24573), .B0(n28610), .B1(n18152), .Y(
        DP_OP_5171J1_127_4278_n81) );
  AOI32XL U22348 ( .A0(n18078), .A1(n24570), .A2(n19693), .B0(n18084), .B1(
        n17936), .Y(DP_OP_5171J1_127_4278_n101) );
  OAI21XL U22349 ( .A0(n19696), .A1(n18154), .B0(n18153), .Y(
        DP_OP_5171J1_127_4278_n90) );
  INVXL U22350 ( .A(affine_2[11]), .Y(DP_OP_5171J1_127_4278_n31) );
  INVXL U22351 ( .A(cs[2]), .Y(n18175) );
  INVXL U22352 ( .A(cs[0]), .Y(n18176) );
  INVXL U22353 ( .A(cs[1]), .Y(n18161) );
  INVXL U22354 ( .A(counter[6]), .Y(n26849) );
  NAND2XL U22355 ( .A(counter[5]), .B(n18773), .Y(n18169) );
  INVXL U22356 ( .A(n18167), .Y(n18168) );
  AOI211XL U22357 ( .A0(n26849), .A1(n18169), .B0(n19242), .C0(n18168), .Y(
        N30145) );
  INVXL U22358 ( .A(n20358), .Y(n18171) );
  AOI211XL U22359 ( .A0(n20600), .A1(n18171), .B0(n19242), .C0(n18773), .Y(
        N30143) );
  INVXL U22360 ( .A(n18187), .Y(n18183) );
  OAI31X2 U22361 ( .A0(n18182), .A1(n18181), .A2(n18180), .B0(n36247), .Y(
        n19180) );
  INVXL U22362 ( .A(ns[1]), .Y(n20616) );
  INVXL U22363 ( .A(n36207), .Y(n36250) );
  NAND2XL U22364 ( .A(n18191), .B(n19006), .Y(n28391) );
  AOI22XL U22365 ( .A0(n22762), .A1(conv_2[389]), .B0(n25299), .B1(conv_2[374]), .Y(n18192) );
  NAND2XL U22366 ( .A(n18193), .B(n18192), .Y(n25618) );
  AOI22XL U22367 ( .A0(n18810), .A1(conv_2[344]), .B0(n16723), .B1(conv_2[359]), .Y(n18195) );
  AOI22XL U22368 ( .A0(n16666), .A1(conv_2[329]), .B0(n22759), .B1(conv_2[314]), .Y(n18194) );
  NAND2XL U22369 ( .A(n18195), .B(n18194), .Y(n25621) );
  NAND2XL U22370 ( .A(N18471), .B(n28290), .Y(n18196) );
  AOI22XL U22371 ( .A0(n21011), .A1(conv_2[209]), .B0(n25299), .B1(conv_2[194]), .Y(n18199) );
  AOI22XL U22372 ( .A0(n16716), .A1(conv_2[224]), .B0(n16723), .B1(conv_2[239]), .Y(n18198) );
  NAND2XL U22373 ( .A(n18199), .B(n18198), .Y(n25628) );
  INVX2 U22374 ( .A(n35196), .Y(n35234) );
  INVXL U22375 ( .A(conv_2[269]), .Y(n28144) );
  INVXL U22376 ( .A(conv_2[254]), .Y(n28153) );
  INVXL U22377 ( .A(N17631), .Y(n19253) );
  AOI22XL U22378 ( .A0(n35269), .A1(n28144), .B0(n28153), .B1(n19253), .Y(
        n25813) );
  AOI222XL U22379 ( .A0(n25813), .A1(n21358), .B0(n16673), .B1(conv_2[299]), 
        .C0(conv_2[284]), .C1(n16716), .Y(n25622) );
  INVXL U22380 ( .A(n25622), .Y(n24778) );
  AOI22XL U22381 ( .A0(n16660), .A1(n25628), .B0(n35234), .B1(n24778), .Y(
        n18212) );
  NOR2X1 U22382 ( .A(n25123), .B(N18014), .Y(n28291) );
  NAND2X2 U22383 ( .A(n28467), .B(n28291), .Y(n35202) );
  INVX4 U22384 ( .A(n35202), .Y(n35181) );
  AOI22XL U22385 ( .A0(n22770), .A1(conv_2[29]), .B0(n22690), .B1(conv_2[14]), 
        .Y(n18201) );
  NAND2XL U22386 ( .A(n18201), .B(n18200), .Y(n25199) );
  INVXL U22387 ( .A(conv_2[89]), .Y(n32677) );
  INVXL U22388 ( .A(conv_2[74]), .Y(n30247) );
  OAI22XL U22389 ( .A0(n19902), .A1(n32677), .B0(n22717), .B1(n30247), .Y(
        n18203) );
  INVXL U22390 ( .A(conv_2[104]), .Y(n30232) );
  INVXL U22391 ( .A(conv_2[119]), .Y(n30254) );
  OAI22XL U22392 ( .A0(n22612), .A1(n30232), .B0(n18321), .B1(n30254), .Y(
        n18202) );
  INVXL U22393 ( .A(conv_2[539]), .Y(n30427) );
  INVXL U22394 ( .A(conv_2[524]), .Y(n29443) );
  AOI22XL U22395 ( .A0(n20735), .A1(n30427), .B0(n29443), .B1(n19253), .Y(
        n25812) );
  INVXL U22396 ( .A(conv_2[509]), .Y(n34016) );
  INVXL U22397 ( .A(conv_2[494]), .Y(n34670) );
  AOI22XL U22398 ( .A0(n35269), .A1(n34016), .B0(n34670), .B1(n18526), .Y(
        n21976) );
  OAI22XL U22399 ( .A0(n25623), .A1(n35239), .B0(n35184), .B1(n25624), .Y(
        n18210) );
  INVXL U22400 ( .A(conv_2[479]), .Y(n27950) );
  INVXL U22401 ( .A(conv_2[464]), .Y(n27964) );
  AOI22XL U22402 ( .A0(n35269), .A1(n27950), .B0(n27964), .B1(n19253), .Y(
        n25819) );
  AOI222XL U22403 ( .A0(n25819), .A1(n36246), .B0(n22759), .B1(conv_2[434]), 
        .C0(n25306), .C1(conv_2[449]), .Y(n25620) );
  INVXL U22404 ( .A(n28290), .Y(n18205) );
  AOI22XL U22405 ( .A0(n22762), .A1(conv_2[149]), .B0(n16723), .B1(conv_2[179]), .Y(n18207) );
  AOI22XL U22406 ( .A0(n16716), .A1(conv_2[164]), .B0(n22690), .B1(conv_2[134]), .Y(n18206) );
  NAND2XL U22407 ( .A(n18207), .B(n18206), .Y(n25619) );
  INVXL U22408 ( .A(n25619), .Y(n25030) );
  NAND2X1 U22409 ( .A(n36245), .B(n23783), .Y(n18208) );
  OAI22XL U22410 ( .A0(n25620), .A1(n35200), .B0(n25030), .B1(n18208), .Y(
        n18209) );
  AOI211XL U22411 ( .A0(n35181), .A1(n25199), .B0(n18210), .C0(n18209), .Y(
        n18211) );
  OAI211XL U22412 ( .A0(n35135), .A1(n24783), .B0(n18212), .C0(n18211), .Y(
        n18449) );
  AOI22XL U22413 ( .A0(n22770), .A1(conv_2[385]), .B0(n16673), .B1(conv_2[415]), .Y(n18213) );
  NAND2XL U22414 ( .A(n18214), .B(n18213), .Y(n25584) );
  AOI22XL U22415 ( .A0(n22762), .A1(conv_2[325]), .B0(n16673), .B1(conv_2[355]), .Y(n18215) );
  NAND2XL U22416 ( .A(n18216), .B(n18215), .Y(n25585) );
  AOI22XL U22417 ( .A0(n36245), .A1(n25584), .B0(n25585), .B1(n26374), .Y(
        n24753) );
  AOI22XL U22418 ( .A0(n20978), .A1(conv_2[85]), .B0(n16662), .B1(conv_2[100]), 
        .Y(n18218) );
  AOI22XL U22419 ( .A0(n25299), .A1(conv_2[70]), .B0(n16673), .B1(conv_2[115]), 
        .Y(n18217) );
  NAND2XL U22420 ( .A(n18218), .B(n18217), .Y(n25588) );
  INVXL U22421 ( .A(conv_2[130]), .Y(n30075) );
  INVXL U22422 ( .A(conv_2[145]), .Y(n30099) );
  INVXL U22423 ( .A(conv_2[175]), .Y(n30897) );
  OAI22XL U22424 ( .A0(n18286), .A1(n30099), .B0(n24039), .B1(n30897), .Y(
        n18219) );
  INVXL U22425 ( .A(n25597), .Y(n24748) );
  AOI22XL U22426 ( .A0(n35195), .A1(n25588), .B0(n35236), .B1(n24748), .Y(
        n18228) );
  INVXL U22427 ( .A(conv_2[430]), .Y(n32894) );
  AOI22XL U22428 ( .A0(n20735), .A1(conv_2[475]), .B0(conv_2[460]), .B1(n18526), .Y(n26038) );
  INVXL U22429 ( .A(conv_2[445]), .Y(n27909) );
  OAI222XL U22430 ( .A0(n32894), .A1(n22717), .B0(n21688), .B1(n26038), .C0(
        n22546), .C1(n27909), .Y(n25183) );
  INVXL U22431 ( .A(conv_2[535]), .Y(n33375) );
  INVXL U22432 ( .A(conv_2[520]), .Y(n27798) );
  INVXL U22433 ( .A(N17631), .Y(n18526) );
  AOI22XL U22434 ( .A0(n20735), .A1(n33375), .B0(n27798), .B1(n18526), .Y(
        n21913) );
  INVXL U22435 ( .A(conv_2[505]), .Y(n36090) );
  INVXL U22436 ( .A(conv_2[490]), .Y(n27751) );
  AOI22XL U22437 ( .A0(n20735), .A1(n36090), .B0(n27751), .B1(n18516), .Y(
        n21914) );
  INVXL U22438 ( .A(conv_2[265]), .Y(n28188) );
  AOI2BB2XL U22439 ( .B0(n20735), .B1(n28188), .A0N(conv_2[250]), .A1N(n35269), 
        .Y(n26032) );
  AOI222XL U22440 ( .A0(n26032), .A1(n21688), .B0(n16673), .B1(conv_2[295]), 
        .C0(conv_2[280]), .C1(n16662), .Y(n25589) );
  OAI22XL U22441 ( .A0(n25586), .A1(n35184), .B0(n25589), .B1(n35196), .Y(
        n18226) );
  INVXL U22442 ( .A(conv_2[205]), .Y(n27858) );
  INVXL U22443 ( .A(conv_2[235]), .Y(n29597) );
  OAI22XL U22444 ( .A0(n19401), .A1(n27858), .B0(n24039), .B1(n29597), .Y(
        n18222) );
  INVXL U22445 ( .A(conv_2[220]), .Y(n30434) );
  INVXL U22446 ( .A(conv_2[190]), .Y(n33459) );
  OAI22XL U22447 ( .A0(n22740), .A1(n30434), .B0(n22717), .B1(n33459), .Y(
        n18221) );
  AOI22XL U22448 ( .A0(n22762), .A1(conv_2[25]), .B0(n16673), .B1(conv_2[55]), 
        .Y(n18224) );
  NAND2XL U22449 ( .A(n18224), .B(n18223), .Y(n25186) );
  INVXL U22450 ( .A(n25186), .Y(n25590) );
  OAI22XL U22451 ( .A0(n25587), .A1(n35198), .B0(n25590), .B1(n35202), .Y(
        n18225) );
  AOI211XL U22452 ( .A0(n16664), .A1(n25183), .B0(n18226), .C0(n18225), .Y(
        n18227) );
  OAI211XL U22453 ( .A0(n35135), .A1(n24753), .B0(n18228), .C0(n18227), .Y(
        n18424) );
  INVXL U22454 ( .A(conv_2[185]), .Y(n29902) );
  INVXL U22455 ( .A(conv_2[200]), .Y(n29945) );
  INVXL U22456 ( .A(conv_2[230]), .Y(n29517) );
  OAI22XL U22457 ( .A0(n22546), .A1(n29945), .B0(n24039), .B1(n29517), .Y(
        n18229) );
  INVX4 U22458 ( .A(n18516), .Y(n20735) );
  INVXL U22459 ( .A(conv_2[470]), .Y(n33896) );
  INVXL U22460 ( .A(conv_2[455]), .Y(n27649) );
  INVXL U22461 ( .A(N17631), .Y(n18634) );
  AOI22XL U22462 ( .A0(n20735), .A1(n33896), .B0(n27649), .B1(n18634), .Y(
        n25897) );
  AOI222XL U22463 ( .A0(n25897), .A1(n36246), .B0(n22759), .B1(conv_2[425]), 
        .C0(n22762), .C1(conv_2[440]), .Y(n25140) );
  INVXL U22464 ( .A(n25140), .Y(n25516) );
  AOI22XL U22465 ( .A0(n20735), .A1(conv_2[530]), .B0(conv_2[515]), .B1(n18634), .Y(n21879) );
  AOI22XL U22466 ( .A0(n20735), .A1(conv_2[500]), .B0(conv_2[485]), .B1(n18634), .Y(n21880) );
  AOI22XL U22467 ( .A0(n16664), .A1(n25516), .B0(n25519), .B1(n35207), .Y(
        n18246) );
  INVXL U22468 ( .A(conv_2[380]), .Y(n29449) );
  INVXL U22469 ( .A(conv_2[365]), .Y(n34568) );
  OAI22XL U22470 ( .A0(n19902), .A1(n29449), .B0(n22717), .B1(n34568), .Y(
        n18232) );
  INVXL U22471 ( .A(conv_2[395]), .Y(n28119) );
  INVXL U22472 ( .A(conv_2[410]), .Y(n33382) );
  OAI22XL U22473 ( .A0(n22740), .A1(n28119), .B0(n24039), .B1(n33382), .Y(
        n18231) );
  AOI22XL U22474 ( .A0(n22762), .A1(conv_2[320]), .B0(n16673), .B1(conv_2[350]), .Y(n18234) );
  NAND2XL U22475 ( .A(n18234), .B(n18233), .Y(n25139) );
  INVXL U22476 ( .A(n25139), .Y(n25512) );
  AOI22XL U22477 ( .A0(n36245), .A1(n25522), .B0(n25512), .B1(n28292), .Y(
        n24735) );
  INVXL U22478 ( .A(conv_2[170]), .Y(n29838) );
  INVXL U22479 ( .A(conv_2[140]), .Y(n34243) );
  INVXL U22480 ( .A(conv_2[125]), .Y(n34128) );
  OAI22XL U22481 ( .A0(n22546), .A1(n34243), .B0(n22717), .B1(n34128), .Y(
        n18235) );
  INVXL U22482 ( .A(conv_2[260]), .Y(n28182) );
  INVXL U22483 ( .A(conv_2[245]), .Y(n28263) );
  AOI22XL U22484 ( .A0(n20735), .A1(n28182), .B0(n28263), .B1(n18634), .Y(
        n25898) );
  AOI222XL U22485 ( .A0(n25898), .A1(n22713), .B0(n16673), .B1(conv_2[290]), 
        .C0(conv_2[275]), .C1(n25289), .Y(n25515) );
  OAI22XL U22486 ( .A0(n25513), .A1(n18208), .B0(n25515), .B1(n35196), .Y(
        n18244) );
  INVXL U22487 ( .A(conv_2[50]), .Y(n27808) );
  INVXL U22488 ( .A(conv_2[20]), .Y(n29080) );
  INVXL U22489 ( .A(conv_2[35]), .Y(n33596) );
  OAI22XL U22490 ( .A0(n22546), .A1(n29080), .B0(n22612), .B1(n33596), .Y(
        n18237) );
  INVXL U22491 ( .A(conv_2[110]), .Y(n28679) );
  INVXL U22492 ( .A(conv_2[80]), .Y(n30183) );
  INVXL U22493 ( .A(conv_2[95]), .Y(n19172) );
  OAI22XL U22494 ( .A0(n22546), .A1(n30183), .B0(n22612), .B1(n19172), .Y(
        n18241) );
  OAI22XL U22495 ( .A0(n25518), .A1(n35202), .B0(n25514), .B1(n35239), .Y(
        n18243) );
  AOI211XL U22496 ( .A0(n28465), .A1(n24735), .B0(n18244), .C0(n18243), .Y(
        n18245) );
  OAI211XL U22497 ( .A0(n25141), .A1(n35198), .B0(n18246), .C0(n18245), .Y(
        n18400) );
  AOI22XL U22498 ( .A0(n22762), .A1(conv_2[79]), .B0(n16673), .B1(conv_2[109]), 
        .Y(n18248) );
  NAND2XL U22499 ( .A(n18248), .B(n18247), .Y(n25135) );
  AOI22XL U22500 ( .A0(n20735), .A1(conv_2[529]), .B0(conv_2[514]), .B1(n18516), .Y(n25936) );
  AOI22XL U22501 ( .A0(n20735), .A1(conv_2[499]), .B0(conv_2[484]), .B1(n18516), .Y(n21866) );
  AOI22XL U22502 ( .A0(n35195), .A1(n25135), .B0(n25501), .B1(n35231), .Y(
        n18263) );
  AOI22XL U22503 ( .A0(n25299), .A1(conv_2[184]), .B0(n16673), .B1(conv_2[229]), .Y(n18250) );
  AOI22XL U22504 ( .A0(n22762), .A1(conv_2[199]), .B0(n16662), .B1(conv_2[214]), .Y(n18249) );
  NAND2XL U22505 ( .A(n18250), .B(n18249), .Y(n25132) );
  INVXL U22506 ( .A(conv_2[259]), .Y(n29413) );
  INVXL U22507 ( .A(conv_2[244]), .Y(n28982) );
  AOI22XL U22508 ( .A0(n20735), .A1(n29413), .B0(n28982), .B1(n18516), .Y(
        n25930) );
  AOI222XL U22509 ( .A0(n25930), .A1(n21688), .B0(n16673), .B1(conv_2[289]), 
        .C0(conv_2[274]), .C1(n25289), .Y(n25502) );
  AOI22XL U22510 ( .A0(n25306), .A1(conv_2[139]), .B0(n22690), .B1(conv_2[124]), .Y(n18251) );
  NAND2XL U22511 ( .A(n18252), .B(n18251), .Y(n25131) );
  INVXL U22512 ( .A(n25131), .Y(n24982) );
  OAI22XL U22513 ( .A0(n25502), .A1(n35196), .B0(n24982), .B1(n18208), .Y(
        n18261) );
  INVXL U22514 ( .A(conv_2[424]), .Y(n29021) );
  AOI22XL U22515 ( .A0(n20735), .A1(conv_2[469]), .B0(conv_2[454]), .B1(n18634), .Y(n21858) );
  INVXL U22516 ( .A(conv_2[439]), .Y(n29033) );
  NAND2XL U22517 ( .A(n16721), .B(n25501), .Y(n25136) );
  AOI22XL U22518 ( .A0(n25306), .A1(conv_2[19]), .B0(n22690), .B1(conv_2[4]), 
        .Y(n18254) );
  NAND2XL U22519 ( .A(n18254), .B(n18253), .Y(n25134) );
  OAI2BB2XL U22520 ( .B0(n26374), .B1(n25136), .A0N(n22362), .A1N(n25134), .Y(
        n18255) );
  AOI21XL U22521 ( .A0(n28292), .A1(n25511), .B0(n18255), .Y(n24727) );
  AOI22XL U22522 ( .A0(n22762), .A1(conv_2[379]), .B0(n16673), .B1(conv_2[409]), .Y(n18257) );
  NAND2XL U22523 ( .A(n18257), .B(n18256), .Y(n25503) );
  AOI22XL U22524 ( .A0(n25299), .A1(conv_2[304]), .B0(n16673), .B1(conv_2[349]), .Y(n18258) );
  NAND2XL U22525 ( .A(n18259), .B(n18258), .Y(n25504) );
  AOI22XL U22526 ( .A0(n36245), .A1(n25503), .B0(n25504), .B1(n26374), .Y(
        n24726) );
  OAI22XL U22527 ( .A0(n24727), .A1(n35159), .B0(n35135), .B1(n24726), .Y(
        n18260) );
  AOI211XL U22528 ( .A0(n16660), .A1(n25132), .B0(n18261), .C0(n18260), .Y(
        n18262) );
  NAND2XL U22529 ( .A(n18263), .B(n18262), .Y(n18451) );
  INVXL U22530 ( .A(conv_2[414]), .Y(n33693) );
  INVXL U22531 ( .A(conv_2[384]), .Y(n28017) );
  INVXL U22532 ( .A(conv_2[399]), .Y(n34640) );
  OAI22XL U22533 ( .A0(n19902), .A1(n28017), .B0(n22612), .B1(n34640), .Y(
        n18264) );
  AOI211XL U22534 ( .A0(n22616), .A1(conv_2[369]), .B0(n18265), .C0(n18264), 
        .Y(n25177) );
  INVXL U22535 ( .A(n25177), .Y(n25570) );
  INVXL U22536 ( .A(conv_2[324]), .Y(n28058) );
  INVXL U22537 ( .A(conv_2[339]), .Y(n35999) );
  OAI22XL U22538 ( .A0(n19902), .A1(n28058), .B0(n22612), .B1(n35999), .Y(
        n18267) );
  INVXL U22539 ( .A(conv_2[309]), .Y(n35972) );
  INVXL U22540 ( .A(conv_2[354]), .Y(n29481) );
  OAI22XL U22541 ( .A0(n22717), .A1(n35972), .B0(n18321), .B1(n29481), .Y(
        n18266) );
  AOI22XL U22542 ( .A0(n20978), .A1(conv_2[144]), .B0(n25299), .B1(conv_2[129]), .Y(n18269) );
  NAND2XL U22543 ( .A(n18269), .B(n18268), .Y(n25175) );
  INVXL U22544 ( .A(conv_2[219]), .Y(n30429) );
  INVXL U22545 ( .A(conv_2[189]), .Y(n29893) );
  OAI22XL U22546 ( .A0(n22740), .A1(n30429), .B0(n22717), .B1(n29893), .Y(
        n18271) );
  INVXL U22547 ( .A(conv_2[204]), .Y(n29932) );
  INVXL U22548 ( .A(conv_2[234]), .Y(n29159) );
  OAI22XL U22549 ( .A0(n19902), .A1(n29932), .B0(n24039), .B1(n29159), .Y(
        n18270) );
  INVXL U22550 ( .A(n25176), .Y(n25571) );
  AOI22XL U22551 ( .A0(n35236), .A1(n25175), .B0(n16660), .B1(n25571), .Y(
        n18279) );
  INVXL U22552 ( .A(conv_2[24]), .Y(n28675) );
  INVXL U22553 ( .A(conv_2[54]), .Y(n28715) );
  OAI22XL U22554 ( .A0(n22546), .A1(n28675), .B0(n24039), .B1(n28715), .Y(
        n18273) );
  INVXL U22555 ( .A(conv_2[39]), .Y(n35864) );
  INVXL U22556 ( .A(conv_2[9]), .Y(n28783) );
  OAI22XL U22557 ( .A0(n22740), .A1(n35864), .B0(n22550), .B1(n28783), .Y(
        n18272) );
  INVXL U22558 ( .A(n25575), .Y(n24061) );
  INVXL U22559 ( .A(conv_2[69]), .Y(n30977) );
  INVXL U22560 ( .A(conv_2[114]), .Y(n30136) );
  OAI22XL U22561 ( .A0(n22717), .A1(n30977), .B0(n24039), .B1(n30136), .Y(
        n18275) );
  INVXL U22562 ( .A(conv_2[84]), .Y(n30174) );
  INVXL U22563 ( .A(conv_2[99]), .Y(n30944) );
  OAI22XL U22564 ( .A0(n19902), .A1(n30174), .B0(n22612), .B1(n30944), .Y(
        n18274) );
  AOI22XL U22565 ( .A0(n20735), .A1(conv_2[534]), .B0(conv_2[519]), .B1(n18526), .Y(n25997) );
  AOI22XL U22566 ( .A0(n20735), .A1(conv_2[504]), .B0(conv_2[489]), .B1(n18526), .Y(n25988) );
  INVXL U22567 ( .A(n25174), .Y(n25577) );
  OAI22XL U22568 ( .A0(n25583), .A1(n35239), .B0(n25577), .B1(n35184), .Y(
        n18277) );
  INVXL U22569 ( .A(conv_2[264]), .Y(n28165) );
  INVXL U22570 ( .A(conv_2[249]), .Y(n33685) );
  AOI22XL U22571 ( .A0(n20735), .A1(n28165), .B0(n33685), .B1(n18516), .Y(
        n20878) );
  AOI222XL U22572 ( .A0(n20878), .A1(n22765), .B0(n16673), .B1(conv_2[294]), 
        .C0(conv_2[279]), .C1(n16662), .Y(n25574) );
  INVXL U22573 ( .A(conv_2[474]), .Y(n30904) );
  INVXL U22574 ( .A(conv_2[459]), .Y(n27654) );
  AOI22XL U22575 ( .A0(n20735), .A1(n30904), .B0(n27654), .B1(n19253), .Y(
        n25992) );
  AOI222XL U22576 ( .A0(n25992), .A1(n36246), .B0(n22759), .B1(conv_2[429]), 
        .C0(n25306), .C1(conv_2[444]), .Y(n25573) );
  OAI22XL U22577 ( .A0(n25574), .A1(n35196), .B0(n25573), .B1(n35200), .Y(
        n18276) );
  AOI211XL U22578 ( .A0(n35181), .A1(n24061), .B0(n18277), .C0(n18276), .Y(
        n18278) );
  OAI211XL U22579 ( .A0(n35135), .A1(n24766), .B0(n18279), .C0(n18278), .Y(
        n18423) );
  NOR4XL U22580 ( .A(n18424), .B(n18400), .C(n18451), .D(n18423), .Y(n18347)
         );
  AOI22XL U22581 ( .A0(n25306), .A1(conv_2[381]), .B0(n16673), .B1(conv_2[411]), .Y(n18280) );
  NAND2XL U22582 ( .A(n18281), .B(n18280), .Y(n25546) );
  AOI22XL U22583 ( .A0(n25306), .A1(conv_2[321]), .B0(n22690), .B1(conv_2[306]), .Y(n18282) );
  NAND2XL U22584 ( .A(n18283), .B(n18282), .Y(n25545) );
  AOI22XL U22585 ( .A0(n36245), .A1(n25546), .B0(n25545), .B1(n28292), .Y(
        n24743) );
  AOI22XL U22586 ( .A0(n25306), .A1(conv_2[141]), .B0(n16673), .B1(conv_2[171]), .Y(n18284) );
  NAND2XL U22587 ( .A(n18285), .B(n18284), .Y(n25547) );
  INVXL U22588 ( .A(conv_2[21]), .Y(n29086) );
  INVXL U22589 ( .A(conv_2[36]), .Y(n27733) );
  INVXL U22590 ( .A(conv_2[6]), .Y(n28777) );
  OAI22XL U22591 ( .A0(n22612), .A1(n27733), .B0(n22717), .B1(n28777), .Y(
        n18287) );
  AOI211XL U22592 ( .A0(n16723), .A1(conv_2[51]), .B0(n18288), .C0(n18287), 
        .Y(n25540) );
  AOI2BB2XL U22593 ( .B0(n35236), .B1(n25547), .A0N(n35202), .A1N(n25540), .Y(
        n18296) );
  AOI22XL U22594 ( .A0(n20735), .A1(conv_2[531]), .B0(conv_2[516]), .B1(n18526), .Y(n25955) );
  AOI22XL U22595 ( .A0(n20735), .A1(conv_2[501]), .B0(conv_2[486]), .B1(n18526), .Y(n25958) );
  AOI22XL U22596 ( .A0(n25306), .A1(conv_2[81]), .B0(n16673), .B1(conv_2[111]), 
        .Y(n18289) );
  NAND2XL U22597 ( .A(n18290), .B(n18289), .Y(n25162) );
  INVXL U22598 ( .A(n25162), .Y(n25550) );
  INVXL U22599 ( .A(conv_2[471]), .Y(n27871) );
  INVXL U22600 ( .A(conv_2[456]), .Y(n30881) );
  AOI22XL U22601 ( .A0(n20735), .A1(n27871), .B0(n30881), .B1(n18634), .Y(
        n25960) );
  AOI222XL U22602 ( .A0(n25960), .A1(n36246), .B0(n22759), .B1(conv_2[426]), 
        .C0(n22770), .C1(conv_2[441]), .Y(n25541) );
  OAI22XL U22603 ( .A0(n25550), .A1(n35239), .B0(n25541), .B1(n35200), .Y(
        n18294) );
  INVXL U22604 ( .A(conv_2[261]), .Y(n34604) );
  INVXL U22605 ( .A(conv_2[246]), .Y(n29148) );
  AOI22XL U22606 ( .A0(n20735), .A1(n34604), .B0(n29148), .B1(n18516), .Y(
        n25949) );
  AOI222XL U22607 ( .A0(n25949), .A1(n22743), .B0(n16673), .B1(conv_2[291]), 
        .C0(conv_2[276]), .C1(n16662), .Y(n25163) );
  INVXL U22608 ( .A(conv_2[231]), .Y(n29178) );
  INVXL U22609 ( .A(conv_2[201]), .Y(n35923) );
  INVXL U22610 ( .A(conv_2[186]), .Y(n29914) );
  OAI22XL U22611 ( .A0(n19902), .A1(n35923), .B0(n22717), .B1(n29914), .Y(
        n18291) );
  OAI22XL U22612 ( .A0(n25163), .A1(n35196), .B0(n25543), .B1(n35198), .Y(
        n18293) );
  AOI211XL U22613 ( .A0(n25542), .A1(n35207), .B0(n18294), .C0(n18293), .Y(
        n18295) );
  OAI211XL U22614 ( .A0(n35135), .A1(n24743), .B0(n18296), .C0(n18295), .Y(
        n18402) );
  AOI22XL U22615 ( .A0(n25306), .A1(conv_2[382]), .B0(n16662), .B1(conv_2[397]), .Y(n18298) );
  AOI22XL U22616 ( .A0(n22690), .A1(conv_2[367]), .B0(n16673), .B1(conv_2[412]), .Y(n18297) );
  NAND2XL U22617 ( .A(n18298), .B(n18297), .Y(n25532) );
  AOI22XL U22618 ( .A0(n22762), .A1(conv_2[322]), .B0(n22690), .B1(conv_2[307]), .Y(n18299) );
  NAND2XL U22619 ( .A(n18300), .B(n18299), .Y(n25533) );
  AOI22XL U22620 ( .A0(n36245), .A1(n25532), .B0(n25533), .B1(n26374), .Y(
        n24738) );
  AOI22XL U22621 ( .A0(n25306), .A1(conv_2[22]), .B0(n25299), .B1(conv_2[7]), 
        .Y(n18301) );
  NAND2XL U22622 ( .A(n18302), .B(n18301), .Y(n25531) );
  AOI22XL U22623 ( .A0(n20735), .A1(conv_2[532]), .B0(conv_2[517]), .B1(n19253), .Y(n25915) );
  AOI22XL U22624 ( .A0(n20735), .A1(conv_2[502]), .B0(conv_2[487]), .B1(n18634), .Y(n20946) );
  AOI22XL U22625 ( .A0(n35181), .A1(n25531), .B0(n25147), .B1(n35207), .Y(
        n18312) );
  AOI22XL U22626 ( .A0(n16666), .A1(conv_2[82]), .B0(n22759), .B1(conv_2[67]), 
        .Y(n18304) );
  NAND2XL U22627 ( .A(n18304), .B(n18303), .Y(n25526) );
  INVXL U22628 ( .A(conv_2[472]), .Y(n27890) );
  INVXL U22629 ( .A(conv_2[457]), .Y(n27670) );
  AOI22XL U22630 ( .A0(n20735), .A1(n27890), .B0(n27670), .B1(n18634), .Y(
        n25918) );
  AOI222XL U22631 ( .A0(n25918), .A1(n36246), .B0(n22690), .B1(conv_2[427]), 
        .C0(n22770), .C1(conv_2[442]), .Y(n25536) );
  OAI22XL U22632 ( .A0(n18526), .A1(conv_2[262]), .B0(conv_2[247]), .B1(n35269), .Y(n20939) );
  INVXL U22633 ( .A(n20939), .Y(n25911) );
  AOI222XL U22634 ( .A0(n25911), .A1(n21688), .B0(n16673), .B1(conv_2[292]), 
        .C0(conv_2[277]), .C1(n25289), .Y(n25527) );
  OAI22XL U22635 ( .A0(n25536), .A1(n35200), .B0(n25527), .B1(n35196), .Y(
        n18310) );
  INVXL U22636 ( .A(conv_2[217]), .Y(n30159) );
  INVXL U22637 ( .A(conv_2[202]), .Y(n29939) );
  INVXL U22638 ( .A(conv_2[187]), .Y(n29890) );
  OAI22XL U22639 ( .A0(n22546), .A1(n29939), .B0(n22717), .B1(n29890), .Y(
        n18305) );
  INVXL U22640 ( .A(conv_2[127]), .Y(n30066) );
  INVXL U22641 ( .A(conv_2[142]), .Y(n35901) );
  INVXL U22642 ( .A(conv_2[157]), .Y(n29867) );
  OAI22XL U22643 ( .A0(n22546), .A1(n35901), .B0(n22612), .B1(n29867), .Y(
        n18307) );
  AOI211XL U22644 ( .A0(n16723), .A1(conv_2[172]), .B0(n18308), .C0(n18307), 
        .Y(n25528) );
  OAI22XL U22645 ( .A0(n25148), .A1(n35198), .B0(n25528), .B1(n18208), .Y(
        n18309) );
  AOI211XL U22646 ( .A0(n35195), .A1(n25526), .B0(n18310), .C0(n18309), .Y(
        n18311) );
  OAI211XL U22647 ( .A0(n35135), .A1(n24738), .B0(n18312), .C0(n18311), .Y(
        n18401) );
  AOI22XL U22648 ( .A0(n22762), .A1(conv_2[383]), .B0(n16673), .B1(conv_2[413]), .Y(n18314) );
  NAND2XL U22649 ( .A(n18314), .B(n18313), .Y(n25561) );
  AOI22XL U22650 ( .A0(n25306), .A1(conv_2[323]), .B0(n22690), .B1(conv_2[308]), .Y(n18316) );
  NAND2XL U22651 ( .A(n18316), .B(n18315), .Y(n25562) );
  AOI22XL U22652 ( .A0(n36245), .A1(n25561), .B0(n25562), .B1(n26374), .Y(
        n24772) );
  AOI22XL U22653 ( .A0(n22762), .A1(conv_2[143]), .B0(n25299), .B1(conv_2[128]), .Y(n18317) );
  NAND2XL U22654 ( .A(n18318), .B(n18317), .Y(n25563) );
  INVXL U22655 ( .A(conv_2[473]), .Y(n27878) );
  INVXL U22656 ( .A(conv_2[458]), .Y(n27676) );
  AOI22XL U22657 ( .A0(n20735), .A1(n27878), .B0(n27676), .B1(n19253), .Y(
        n25976) );
  AOI222XL U22658 ( .A0(n25976), .A1(n36246), .B0(n18658), .B1(conv_2[428]), 
        .C0(n22770), .C1(conv_2[443]), .Y(n25557) );
  INVXL U22659 ( .A(n25557), .Y(n25010) );
  AOI22XL U22660 ( .A0(n35236), .A1(n25563), .B0(n16664), .B1(n25010), .Y(
        n18329) );
  AOI22XL U22661 ( .A0(n22762), .A1(conv_2[23]), .B0(n16673), .B1(conv_2[53]), 
        .Y(n18320) );
  NAND2XL U22662 ( .A(n18320), .B(n18319), .Y(n25558) );
  INVXL U22663 ( .A(conv_2[233]), .Y(n29188) );
  INVXL U22664 ( .A(conv_2[203]), .Y(n35930) );
  INVXL U22665 ( .A(conv_2[188]), .Y(n35916) );
  OAI22XL U22666 ( .A0(n22546), .A1(n35930), .B0(n22717), .B1(n35916), .Y(
        n18322) );
  INVXL U22667 ( .A(conv_2[68]), .Y(n30111) );
  INVXL U22668 ( .A(conv_2[113]), .Y(n35893) );
  OAI22XL U22669 ( .A0(n22717), .A1(n30111), .B0(n24039), .B1(n35893), .Y(
        n18325) );
  INVXL U22670 ( .A(conv_2[83]), .Y(n35878) );
  INVXL U22671 ( .A(conv_2[98]), .Y(n30224) );
  OAI22XL U22672 ( .A0(n19902), .A1(n35878), .B0(n22612), .B1(n30224), .Y(
        n18324) );
  OAI22XL U22673 ( .A0(n25566), .A1(n35198), .B0(n25556), .B1(n35239), .Y(
        n18327) );
  INVXL U22674 ( .A(conv_2[263]), .Y(n28195) );
  INVXL U22675 ( .A(conv_2[248]), .Y(n29154) );
  AOI22XL U22676 ( .A0(n20735), .A1(n28195), .B0(n29154), .B1(n19253), .Y(
        n25969) );
  AOI222XL U22677 ( .A0(n25969), .A1(n22765), .B0(n16673), .B1(conv_2[293]), 
        .C0(conv_2[278]), .C1(n25289), .Y(n25559) );
  AOI22XL U22678 ( .A0(n20735), .A1(conv_2[533]), .B0(conv_2[518]), .B1(n18526), .Y(n20803) );
  AOI22XL U22679 ( .A0(n20735), .A1(conv_2[503]), .B0(conv_2[488]), .B1(n18634), .Y(n21931) );
  INVXL U22680 ( .A(n25560), .Y(n24767) );
  OAI22XL U22681 ( .A0(n25559), .A1(n35196), .B0(n24767), .B1(n35184), .Y(
        n18326) );
  AOI211XL U22682 ( .A0(n35181), .A1(n25558), .B0(n18327), .C0(n18326), .Y(
        n18328) );
  OAI211XL U22683 ( .A0(n35135), .A1(n24772), .B0(n18329), .C0(n18328), .Y(
        n18442) );
  AOI22XL U22684 ( .A0(n22762), .A1(conv_2[386]), .B0(n16673), .B1(conv_2[416]), .Y(n18331) );
  NAND2XL U22685 ( .A(n18331), .B(n18330), .Y(n25004) );
  AOI22XL U22686 ( .A0(n22762), .A1(conv_2[326]), .B0(n16673), .B1(conv_2[356]), .Y(n18332) );
  NAND2XL U22687 ( .A(n18333), .B(n18332), .Y(n25599) );
  AOI22XL U22688 ( .A0(n36245), .A1(n25004), .B0(n25599), .B1(n28292), .Y(
        n24761) );
  AOI22XL U22689 ( .A0(n22762), .A1(conv_2[86]), .B0(n16673), .B1(conv_2[116]), 
        .Y(n18334) );
  NAND2XL U22690 ( .A(n18335), .B(n18334), .Y(n25601) );
  INVXL U22691 ( .A(conv_2[476]), .Y(n27896) );
  INVXL U22692 ( .A(conv_2[461]), .Y(n27659) );
  AOI22XL U22693 ( .A0(n20735), .A1(n27896), .B0(n27659), .B1(n18516), .Y(
        n26011) );
  AOI222XL U22694 ( .A0(n26011), .A1(n36246), .B0(n22759), .B1(conv_2[431]), 
        .C0(n25306), .C1(conv_2[446]), .Y(n25154) );
  INVXL U22695 ( .A(n25154), .Y(n25598) );
  AOI22XL U22696 ( .A0(n35195), .A1(n25601), .B0(n16664), .B1(n25598), .Y(
        n18345) );
  AOI22XL U22697 ( .A0(n25299), .A1(conv_2[131]), .B0(n16673), .B1(conv_2[176]), .Y(n18337) );
  AOI22XL U22698 ( .A0(n22762), .A1(conv_2[146]), .B0(n16662), .B1(conv_2[161]), .Y(n18336) );
  NAND2XL U22699 ( .A(n18337), .B(n18336), .Y(n25600) );
  INVXL U22700 ( .A(conv_2[191]), .Y(n29908) );
  INVXL U22701 ( .A(conv_2[221]), .Y(n30437) );
  INVXL U22702 ( .A(conv_2[236]), .Y(n30936) );
  OAI22XL U22703 ( .A0(n22612), .A1(n30437), .B0(n24039), .B1(n30936), .Y(
        n18338) );
  AOI211XL U22704 ( .A0(n25306), .A1(conv_2[206]), .B0(n18339), .C0(n18338), 
        .Y(n25603) );
  AOI22XL U22705 ( .A0(n20735), .A1(conv_2[536]), .B0(conv_2[521]), .B1(n18526), .Y(n26027) );
  AOI22XL U22706 ( .A0(n20735), .A1(conv_2[506]), .B0(conv_2[491]), .B1(n19253), .Y(n26009) );
  INVXL U22707 ( .A(n25156), .Y(n25602) );
  OAI22XL U22708 ( .A0(n25603), .A1(n35198), .B0(n25602), .B1(n35184), .Y(
        n18343) );
  INVXL U22709 ( .A(conv_2[266]), .Y(n28171) );
  INVXL U22710 ( .A(conv_2[251]), .Y(n35944) );
  AOI22XL U22711 ( .A0(n20735), .A1(n28171), .B0(n35944), .B1(n19253), .Y(
        n26007) );
  AOI222XL U22712 ( .A0(n26007), .A1(n22765), .B0(n16673), .B1(conv_2[296]), 
        .C0(conv_2[281]), .C1(n16662), .Y(n25155) );
  INVXL U22713 ( .A(conv_2[41]), .Y(n29622) );
  INVXL U22714 ( .A(conv_2[56]), .Y(n30161) );
  OAI22XL U22715 ( .A0(n22740), .A1(n29622), .B0(n24039), .B1(n30161), .Y(
        n18341) );
  INVXL U22716 ( .A(conv_2[26]), .Y(n27841) );
  INVXL U22717 ( .A(conv_2[11]), .Y(n27696) );
  OAI22XL U22718 ( .A0(n22546), .A1(n27841), .B0(n22550), .B1(n27696), .Y(
        n18340) );
  OAI22XL U22719 ( .A0(n25155), .A1(n35196), .B0(n25604), .B1(n35202), .Y(
        n18342) );
  AOI211XL U22720 ( .A0(n35236), .A1(n25600), .B0(n18343), .C0(n18342), .Y(
        n18344) );
  OAI211XL U22721 ( .A0(n35135), .A1(n24761), .B0(n18345), .C0(n18344), .Y(
        n18425) );
  NOR4XL U22722 ( .A(n18402), .B(n18401), .C(n18442), .D(n18425), .Y(n18346)
         );
  AOI21XL U22723 ( .A0(n18347), .A1(n18346), .B0(pool[89]), .Y(n18405) );
  AOI22XL U22724 ( .A0(n20735), .A1(conv_2[528]), .B0(conv_2[513]), .B1(n18516), .Y(n21818) );
  AOI22XL U22725 ( .A0(n20735), .A1(conv_2[498]), .B0(conv_2[483]), .B1(n18516), .Y(n25836) );
  NAND2XL U22726 ( .A(n16721), .B(n24956), .Y(n25109) );
  AOI22XL U22727 ( .A0(n16662), .A1(conv_2[33]), .B0(n16673), .B1(conv_2[48]), 
        .Y(n18349) );
  NAND2XL U22728 ( .A(n18349), .B(n18348), .Y(n25107) );
  INVXL U22729 ( .A(conv_2[423]), .Y(n32874) );
  AOI22XL U22730 ( .A0(n35269), .A1(conv_2[468]), .B0(conv_2[453]), .B1(n18526), .Y(n21819) );
  INVXL U22731 ( .A(conv_2[438]), .Y(n29558) );
  OAI222XL U22732 ( .A0(n32874), .A1(n22717), .B0(n22743), .B1(n21819), .C0(
        n22546), .C1(n29558), .Y(n25469) );
  AOI22XL U22733 ( .A0(n22362), .A1(n25107), .B0(n26374), .B1(n25469), .Y(
        n18350) );
  AOI22XL U22734 ( .A0(n22762), .A1(conv_2[378]), .B0(n16662), .B1(conv_2[393]), .Y(n18352) );
  AOI22XL U22735 ( .A0(n25299), .A1(conv_2[363]), .B0(n16673), .B1(conv_2[408]), .Y(n18351) );
  NAND2XL U22736 ( .A(n18352), .B(n18351), .Y(n25467) );
  AOI22XL U22737 ( .A0(n16662), .A1(conv_2[333]), .B0(n22690), .B1(conv_2[303]), .Y(n18354) );
  NAND2XL U22738 ( .A(n18354), .B(n18353), .Y(n25468) );
  AOI22XL U22739 ( .A0(n36245), .A1(n25467), .B0(n25468), .B1(n28292), .Y(
        n24704) );
  AOI22XL U22740 ( .A0(n16662), .A1(conv_2[153]), .B0(n22690), .B1(conv_2[123]), .Y(n18356) );
  NAND2XL U22741 ( .A(n18356), .B(n18355), .Y(n25104) );
  INVXL U22742 ( .A(conv_2[258]), .Y(n32987) );
  INVXL U22743 ( .A(conv_2[243]), .Y(n23161) );
  AOI22XL U22744 ( .A0(n35269), .A1(n32987), .B0(n23161), .B1(n18634), .Y(
        n25838) );
  AOI222XL U22745 ( .A0(n25838), .A1(n21688), .B0(n18810), .B1(conv_2[273]), 
        .C0(conv_2[288]), .C1(n16673), .Y(n24959) );
  INVXL U22746 ( .A(n24959), .Y(n25470) );
  AOI22XL U22747 ( .A0(n35236), .A1(n25104), .B0(n35234), .B1(n25470), .Y(
        n18362) );
  AOI22XL U22748 ( .A0(n16662), .A1(conv_2[93]), .B0(n22759), .B1(conv_2[63]), 
        .Y(n18358) );
  AOI22XL U22749 ( .A0(n22762), .A1(conv_2[78]), .B0(n16673), .B1(conv_2[108]), 
        .Y(n18357) );
  NAND2XL U22750 ( .A(n18358), .B(n18357), .Y(n25108) );
  AOI22XL U22751 ( .A0(n22762), .A1(conv_2[198]), .B0(n16662), .B1(conv_2[213]), .Y(n18360) );
  AOI22XL U22752 ( .A0(n25299), .A1(conv_2[183]), .B0(n16673), .B1(conv_2[228]), .Y(n18359) );
  NAND2XL U22753 ( .A(n18360), .B(n18359), .Y(n25105) );
  AOI22XL U22754 ( .A0(n35195), .A1(n25108), .B0(n18197), .B1(n25105), .Y(
        n18361) );
  OAI211XL U22755 ( .A0(n24962), .A1(n35143), .B0(n18362), .C0(n18361), .Y(
        n18363) );
  INVXL U22756 ( .A(pool[87]), .Y(n34941) );
  INVXL U22757 ( .A(conv_2[527]), .Y(n27057) );
  AOI2BB2XL U22758 ( .B0(n20735), .B1(n27057), .A0N(conv_2[512]), .A1N(n35269), 
        .Y(n20981) );
  INVXL U22759 ( .A(conv_2[497]), .Y(n30323) );
  INVXL U22760 ( .A(conv_2[482]), .Y(n30342) );
  AOI22XL U22761 ( .A0(n20735), .A1(n30323), .B0(n30342), .B1(n18634), .Y(
        n25854) );
  AOI22XL U22762 ( .A0(n22762), .A1(conv_2[137]), .B0(n22690), .B1(conv_2[122]), .Y(n18365) );
  NAND2XL U22763 ( .A(n18366), .B(n18365), .Y(n25122) );
  AOI22XL U22764 ( .A0(n25299), .A1(conv_2[182]), .B0(n16673), .B1(conv_2[227]), .Y(n18367) );
  NAND2XL U22765 ( .A(n18368), .B(n18367), .Y(n24715) );
  AOI22XL U22766 ( .A0(n35236), .A1(n25122), .B0(n16660), .B1(n24715), .Y(
        n18381) );
  INVXL U22767 ( .A(conv_2[257]), .Y(n27049) );
  AOI2BB2X1 U22768 ( .B0(n20735), .B1(n27049), .A0N(conv_2[242]), .A1N(n35269), 
        .Y(n25867) );
  AOI222XL U22769 ( .A0(n25867), .A1(n22713), .B0(n18810), .B1(conv_2[272]), 
        .C0(conv_2[287]), .C1(n16673), .Y(n25491) );
  AOI22XL U22770 ( .A0(n22762), .A1(conv_2[77]), .B0(n16673), .B1(conv_2[107]), 
        .Y(n18369) );
  OAI22XL U22771 ( .A0(n25491), .A1(n35196), .B0(n25124), .B1(n35239), .Y(
        n18379) );
  AOI22XL U22772 ( .A0(n25299), .A1(conv_2[2]), .B0(n16673), .B1(conv_2[47]), 
        .Y(n18372) );
  NAND2XL U22773 ( .A(n18372), .B(n18371), .Y(n25127) );
  INVXL U22774 ( .A(conv_2[467]), .Y(n30336) );
  INVXL U22775 ( .A(conv_2[452]), .Y(n30017) );
  AOI22XL U22776 ( .A0(n35269), .A1(n30336), .B0(n30017), .B1(n18526), .Y(
        n25855) );
  AOI222XL U22777 ( .A0(n25855), .A1(n36246), .B0(n22690), .B1(conv_2[422]), 
        .C0(n22770), .C1(conv_2[437]), .Y(n25490) );
  INVXL U22778 ( .A(n25490), .Y(n18373) );
  NOR2XL U22779 ( .A(N18014), .B(n18815), .Y(n28289) );
  AOI222XL U22780 ( .A0(n25127), .A1(n28291), .B0(n18373), .B1(n28290), .C0(
        n25496), .C1(n28289), .Y(n24717) );
  AOI22XL U22781 ( .A0(n16662), .A1(conv_2[392]), .B0(n22690), .B1(conv_2[362]), .Y(n18375) );
  AOI22XL U22782 ( .A0(n22762), .A1(conv_2[377]), .B0(n16673), .B1(conv_2[407]), .Y(n18374) );
  NAND2XL U22783 ( .A(n18375), .B(n18374), .Y(n25488) );
  AOI22XL U22784 ( .A0(n16662), .A1(conv_2[332]), .B0(n16673), .B1(conv_2[347]), .Y(n18376) );
  NAND2XL U22785 ( .A(n18377), .B(n18376), .Y(n25489) );
  AOI22XL U22786 ( .A0(n36245), .A1(n25488), .B0(n25489), .B1(n26374), .Y(
        n24716) );
  OAI22XL U22787 ( .A0(N18471), .A1(n24717), .B0(n24716), .B1(n35135), .Y(
        n18378) );
  OAI211XL U22788 ( .A0(n25119), .A1(n35143), .B0(n18381), .C0(n18380), .Y(
        n34939) );
  AOI22XL U22789 ( .A0(n22762), .A1(conv_2[16]), .B0(n22616), .B1(conv_2[1]), 
        .Y(n18383) );
  NAND2XL U22790 ( .A(n18383), .B(n18382), .Y(n24972) );
  INVXL U22791 ( .A(conv_2[526]), .Y(n29780) );
  INVXL U22792 ( .A(conv_2[511]), .Y(n29804) );
  AOI22XL U22793 ( .A0(n20735), .A1(n29780), .B0(n29804), .B1(n19253), .Y(
        n25874) );
  INVXL U22794 ( .A(conv_2[496]), .Y(n34237) );
  INVXL U22795 ( .A(conv_2[481]), .Y(n30293) );
  AOI22XL U22796 ( .A0(n20735), .A1(n34237), .B0(n30293), .B1(n18634), .Y(
        n21849) );
  AOI21XL U22797 ( .A0(n36244), .A1(n24972), .B0(n25116), .Y(n25112) );
  INVXL U22798 ( .A(conv_2[466]), .Y(n30297) );
  INVXL U22799 ( .A(conv_2[451]), .Y(n29792) );
  OAI22XL U22800 ( .A0(n19253), .A1(n30297), .B0(n29792), .B1(n35269), .Y(
        n25876) );
  AOI222XL U22801 ( .A0(conv_2[421]), .A1(n18658), .B0(n36246), .B1(n25876), 
        .C0(n22770), .C1(conv_2[436]), .Y(n25477) );
  AOI22XL U22802 ( .A0(n36245), .A1(n25112), .B0(n25477), .B1(n26374), .Y(
        n24714) );
  AOI22XL U22803 ( .A0(n16666), .A1(conv_2[76]), .B0(n16662), .B1(conv_2[91]), 
        .Y(n18385) );
  AOI22XL U22804 ( .A0(n18658), .A1(conv_2[61]), .B0(n16673), .B1(conv_2[106]), 
        .Y(n18384) );
  NAND2XL U22805 ( .A(n18385), .B(n18384), .Y(n24709) );
  OAI22XL U22806 ( .A0(n24971), .A1(n35143), .B0(n25113), .B1(n35239), .Y(
        n18397) );
  AOI22XL U22807 ( .A0(n22616), .A1(conv_2[361]), .B0(n16673), .B1(conv_2[406]), .Y(n18387) );
  NAND2XL U22808 ( .A(n18387), .B(n18386), .Y(n25478) );
  AOI22XL U22809 ( .A0(n22762), .A1(conv_2[316]), .B0(n16662), .B1(conv_2[331]), .Y(n18389) );
  AOI22XL U22810 ( .A0(n22616), .A1(conv_2[301]), .B0(n16673), .B1(conv_2[346]), .Y(n18388) );
  NAND2XL U22811 ( .A(n18389), .B(n18388), .Y(n25479) );
  AOI22XL U22812 ( .A0(n36245), .A1(n25478), .B0(n25479), .B1(n28292), .Y(
        n24708) );
  AOI22XL U22813 ( .A0(n22762), .A1(conv_2[136]), .B0(n16673), .B1(conv_2[166]), .Y(n18391) );
  NAND2XL U22814 ( .A(n18391), .B(n18390), .Y(n25114) );
  INVXL U22815 ( .A(conv_2[271]), .Y(n24554) );
  AOI22XL U22816 ( .A0(n20735), .A1(conv_2[256]), .B0(conv_2[241]), .B1(n19253), .Y(n25873) );
  INVXL U22817 ( .A(conv_2[286]), .Y(n30305) );
  AOI22XL U22818 ( .A0(n35236), .A1(n25114), .B0(n35234), .B1(n25487), .Y(
        n18395) );
  AOI22XL U22819 ( .A0(n22762), .A1(conv_2[196]), .B0(n18658), .B1(conv_2[181]), .Y(n18393) );
  NAND2XL U22820 ( .A(n18393), .B(n18392), .Y(n25115) );
  NAND2XL U22821 ( .A(n16660), .B(n25115), .Y(n18394) );
  OAI211XL U22822 ( .A0(n24708), .A1(n35135), .B0(n18395), .C0(n18394), .Y(
        n18396) );
  AOI222XL U22823 ( .A0(pool[85]), .A1(pool[86]), .B0(pool[85]), .B1(n22200), 
        .C0(pool[86]), .C1(n22200), .Y(n18398) );
  AOI222XL U22824 ( .A0(n34941), .A1(n34939), .B0(n34941), .B1(n18398), .C0(
        n34939), .C1(n18398), .Y(n18399) );
  AOI222XL U22825 ( .A0(n34942), .A1(pool[88]), .B0(n34942), .B1(n18399), .C0(
        pool[88]), .C1(n18399), .Y(n18404) );
  NAND4XL U22826 ( .A(n18402), .B(n18401), .C(n18400), .D(n18451), .Y(n18403)
         );
  INVXL U22827 ( .A(conv_2[433]), .Y(n28916) );
  AOI22XL U22828 ( .A0(n35269), .A1(conv_2[478]), .B0(conv_2[463]), .B1(n19253), .Y(n26087) );
  INVXL U22829 ( .A(conv_2[448]), .Y(n34734) );
  OAI222XL U22830 ( .A0(n28916), .A1(n22717), .B0(n21358), .B1(n26087), .C0(
        n19401), .C1(n34734), .Y(n25647) );
  INVXL U22831 ( .A(conv_2[223]), .Y(n33267) );
  INVXL U22832 ( .A(conv_2[193]), .Y(n29952) );
  INVXL U22833 ( .A(conv_2[238]), .Y(n33094) );
  OAI22XL U22834 ( .A0(n22717), .A1(n29952), .B0(n18321), .B1(n33094), .Y(
        n18406) );
  AOI211XL U22835 ( .A0(conv_2[208]), .A1(n16666), .B0(n18407), .C0(n18406), 
        .Y(n25654) );
  INVXL U22836 ( .A(conv_2[538]), .Y(n30421) );
  INVXL U22837 ( .A(conv_2[523]), .Y(n29437) );
  AOI22XL U22838 ( .A0(n20735), .A1(n30421), .B0(n29437), .B1(n19253), .Y(
        n21059) );
  INVXL U22839 ( .A(conv_2[508]), .Y(n34010) );
  INVXL U22840 ( .A(conv_2[493]), .Y(n34662) );
  AOI22XL U22841 ( .A0(n20735), .A1(n34010), .B0(n34662), .B1(n18516), .Y(
        n22012) );
  OAI22XL U22842 ( .A0(n25654), .A1(n35198), .B0(n25652), .B1(n35184), .Y(
        n18421) );
  AOI22XL U22843 ( .A0(n25299), .A1(conv_2[373]), .B0(n16673), .B1(conv_2[418]), .Y(n18409) );
  AOI22XL U22844 ( .A0(n22762), .A1(conv_2[388]), .B0(n16662), .B1(conv_2[403]), .Y(n18408) );
  NAND2XL U22845 ( .A(n18409), .B(n18408), .Y(n25649) );
  INVXL U22846 ( .A(conv_2[343]), .Y(n34221) );
  INVXL U22847 ( .A(conv_2[328]), .Y(n33231) );
  INVXL U22848 ( .A(conv_2[358]), .Y(n29478) );
  OAI22XL U22849 ( .A0(n18286), .A1(n33231), .B0(n18321), .B1(n29478), .Y(
        n18410) );
  AOI211XL U22850 ( .A0(n22759), .A1(conv_2[313]), .B0(n18411), .C0(n18410), 
        .Y(n25653) );
  AOI22XL U22851 ( .A0(n16662), .A1(conv_2[43]), .B0(n16673), .B1(conv_2[58]), 
        .Y(n18413) );
  AOI22XL U22852 ( .A0(n16666), .A1(conv_2[28]), .B0(n22690), .B1(conv_2[13]), 
        .Y(n18412) );
  NAND2XL U22853 ( .A(n18413), .B(n18412), .Y(n25651) );
  AOI22XL U22854 ( .A0(n22762), .A1(conv_2[148]), .B0(n16673), .B1(conv_2[178]), .Y(n18415) );
  AOI22XL U22855 ( .A0(n16662), .A1(conv_2[163]), .B0(n25299), .B1(conv_2[133]), .Y(n18414) );
  NAND2XL U22856 ( .A(n18415), .B(n18414), .Y(n25648) );
  AOI22XL U22857 ( .A0(n35181), .A1(n25651), .B0(n35236), .B1(n25648), .Y(
        n18419) );
  AOI22XL U22858 ( .A0(n25299), .A1(conv_2[73]), .B0(n16673), .B1(conv_2[118]), 
        .Y(n18417) );
  NAND2XL U22859 ( .A(n18417), .B(n18416), .Y(n25657) );
  INVXL U22860 ( .A(conv_2[268]), .Y(n28201) );
  INVXL U22861 ( .A(conv_2[253]), .Y(n34148) );
  AOI22XL U22862 ( .A0(n20735), .A1(n28201), .B0(n34148), .B1(n19253), .Y(
        n26080) );
  AOI222XL U22863 ( .A0(n26080), .A1(n22743), .B0(n16673), .B1(conv_2[298]), 
        .C0(conv_2[283]), .C1(n25289), .Y(n25211) );
  INVXL U22864 ( .A(n25211), .Y(n25650) );
  AOI22XL U22865 ( .A0(n35195), .A1(n25657), .B0(n35234), .B1(n25650), .Y(
        n18418) );
  OAI211XL U22866 ( .A0(n35135), .A1(n24793), .B0(n18419), .C0(n18418), .Y(
        n18420) );
  AOI211XL U22867 ( .A0(n16664), .A1(n25647), .B0(n18421), .C0(n18420), .Y(
        n18422) );
  INVXL U22868 ( .A(n18422), .Y(n18444) );
  INVXL U22869 ( .A(conv_2[87]), .Y(n30926) );
  INVXL U22870 ( .A(conv_2[117]), .Y(n34368) );
  OAI22XL U22871 ( .A0(n19902), .A1(n30926), .B0(n18321), .B1(n34368), .Y(
        n18427) );
  INVXL U22872 ( .A(conv_2[102]), .Y(n30228) );
  INVXL U22873 ( .A(conv_2[72]), .Y(n33737) );
  OAI22XL U22874 ( .A0(n22612), .A1(n30228), .B0(n22550), .B1(n33737), .Y(
        n18426) );
  AOI22XL U22875 ( .A0(n16716), .A1(conv_2[42]), .B0(n25299), .B1(conv_2[12]), 
        .Y(n18429) );
  AOI22XL U22876 ( .A0(n21011), .A1(conv_2[27]), .B0(n16673), .B1(conv_2[57]), 
        .Y(n18428) );
  NAND2XL U22877 ( .A(n18429), .B(n18428), .Y(n25643) );
  AOI22XL U22878 ( .A0(n25299), .A1(conv_2[192]), .B0(n16673), .B1(conv_2[237]), .Y(n18431) );
  AOI22XL U22879 ( .A0(n22770), .A1(conv_2[207]), .B0(n16662), .B1(conv_2[222]), .Y(n18430) );
  NAND2XL U22880 ( .A(n18431), .B(n18430), .Y(n25632) );
  AOI22XL U22881 ( .A0(n35181), .A1(n25643), .B0(n16660), .B1(n25632), .Y(
        n18441) );
  AOI22XL U22882 ( .A0(n22762), .A1(conv_2[387]), .B0(n22759), .B1(conv_2[372]), .Y(n18433) );
  AOI22XL U22883 ( .A0(n16662), .A1(conv_2[402]), .B0(n16673), .B1(conv_2[417]), .Y(n18432) );
  NAND2XL U22884 ( .A(n18433), .B(n18432), .Y(n25638) );
  AOI22XL U22885 ( .A0(n16662), .A1(conv_2[342]), .B0(n22690), .B1(conv_2[312]), .Y(n18435) );
  AOI22XL U22886 ( .A0(n25306), .A1(conv_2[327]), .B0(n16673), .B1(conv_2[357]), .Y(n18434) );
  NAND2XL U22887 ( .A(n18435), .B(n18434), .Y(n25639) );
  OAI22XL U22888 ( .A0(n26374), .A1(n25638), .B0(n25639), .B1(n36245), .Y(
        n24788) );
  INVXL U22889 ( .A(n24788), .Y(n24122) );
  INVXL U22890 ( .A(conv_2[537]), .Y(n28253) );
  INVXL U22891 ( .A(conv_2[522]), .Y(n28203) );
  AOI22XL U22892 ( .A0(n35269), .A1(n28253), .B0(n28203), .B1(n18516), .Y(
        n21997) );
  INVXL U22893 ( .A(conv_2[507]), .Y(n33173) );
  INVXL U22894 ( .A(conv_2[492]), .Y(n34131) );
  AOI22XL U22895 ( .A0(n35269), .A1(n33173), .B0(n34131), .B1(n19253), .Y(
        n26065) );
  INVXL U22896 ( .A(conv_2[477]), .Y(n27946) );
  INVXL U22897 ( .A(conv_2[462]), .Y(n27679) );
  AOI22XL U22898 ( .A0(n20735), .A1(n27946), .B0(n27679), .B1(n18516), .Y(
        n26067) );
  AOI222XL U22899 ( .A0(n26067), .A1(n36246), .B0(n22759), .B1(conv_2[432]), 
        .C0(n25306), .C1(conv_2[447]), .Y(n25634) );
  OAI22XL U22900 ( .A0(n25636), .A1(n35184), .B0(n25634), .B1(n35200), .Y(
        n18439) );
  INVXL U22901 ( .A(conv_2[267]), .Y(n28176) );
  INVXL U22902 ( .A(conv_2[252]), .Y(n29460) );
  AOI22XL U22903 ( .A0(n35269), .A1(n28176), .B0(n29460), .B1(n18516), .Y(
        n26064) );
  AOI222XL U22904 ( .A0(n26064), .A1(n21358), .B0(n16673), .B1(conv_2[297]), 
        .C0(conv_2[282]), .C1(n16662), .Y(n25637) );
  AOI22XL U22905 ( .A0(n25299), .A1(conv_2[132]), .B0(n16673), .B1(conv_2[177]), .Y(n18437) );
  AOI22XL U22906 ( .A0(n22762), .A1(conv_2[147]), .B0(n16716), .B1(conv_2[162]), .Y(n18436) );
  NAND2XL U22907 ( .A(n18437), .B(n18436), .Y(n25635) );
  INVXL U22908 ( .A(n25635), .Y(n24125) );
  OAI22XL U22909 ( .A0(n25637), .A1(n35196), .B0(n24125), .B1(n18208), .Y(
        n18438) );
  AOI211XL U22910 ( .A0(n28465), .A1(n24122), .B0(n18439), .C0(n18438), .Y(
        n18440) );
  OAI211XL U22911 ( .A0(n25205), .A1(n35239), .B0(n18441), .C0(n18440), .Y(
        n18445) );
  NAND4XL U22912 ( .A(pool[89]), .B(n18443), .C(n18445), .D(n18442), .Y(n18447) );
  NOR3XL U22913 ( .A(pool[89]), .B(n18445), .C(n18444), .Y(n18446) );
  OAI22XL U22914 ( .A0(n34940), .A1(n18451), .B0(pool[89]), .B1(n34943), .Y(
        n18452) );
  INVXL U22915 ( .A(n18452), .Y(N29305) );
  NAND2XL U22916 ( .A(n26207), .B(n20755), .Y(n28571) );
  INVXL U22917 ( .A(n28571), .Y(n28551) );
  AOI22XL U22918 ( .A0(n20735), .A1(conv_3[530]), .B0(conv_3[515]), .B1(n18634), .Y(n21242) );
  AOI22XL U22919 ( .A0(n20735), .A1(conv_3[500]), .B0(conv_3[485]), .B1(n18516), .Y(n21236) );
  INVXL U22920 ( .A(n35045), .Y(n28309) );
  INVXL U22921 ( .A(conv_3[260]), .Y(n29117) );
  INVXL U22922 ( .A(conv_3[245]), .Y(n34249) );
  AOI22XL U22923 ( .A0(n20735), .A1(n29117), .B0(n34249), .B1(n18516), .Y(
        n21235) );
  AOI222XL U22924 ( .A0(n21235), .A1(n21688), .B0(n16673), .B1(conv_3[290]), 
        .C0(conv_3[275]), .C1(n25289), .Y(n26190) );
  OAI22XL U22925 ( .A0(n28551), .A1(n28309), .B0(n26190), .B1(n34981), .Y(
        n18470) );
  OAI22XL U22926 ( .A0(n18634), .A1(conv_3[470]), .B0(conv_3[455]), .B1(n35269), .Y(n21238) );
  INVXL U22927 ( .A(n21238), .Y(n20503) );
  AOI222XL U22928 ( .A0(n20503), .A1(n36246), .B0(n22759), .B1(conv_3[425]), 
        .C0(n22762), .C1(conv_3[440]), .Y(n25748) );
  INVXL U22929 ( .A(n26263), .Y(n34958) );
  INVX2 U22930 ( .A(n16668), .Y(n22690) );
  AOI22XL U22931 ( .A0(n16662), .A1(conv_3[35]), .B0(n22690), .B1(conv_3[5]), 
        .Y(n18453) );
  NAND2XL U22932 ( .A(n18454), .B(n18453), .Y(n26193) );
  INVXL U22933 ( .A(n26193), .Y(n35042) );
  OAI22XL U22934 ( .A0(n25748), .A1(n34958), .B0(n35042), .B1(n35198), .Y(
        n18469) );
  INVXL U22935 ( .A(conv_3[155]), .Y(n32289) );
  INVXL U22936 ( .A(conv_3[125]), .Y(n31403) );
  OAI22XL U22937 ( .A0(n22740), .A1(n32289), .B0(n22717), .B1(n31403), .Y(
        n18456) );
  INVXL U22938 ( .A(conv_3[140]), .Y(n34400) );
  INVXL U22939 ( .A(conv_3[170]), .Y(n31589) );
  OAI22XL U22940 ( .A0(n19902), .A1(n34400), .B0(n18321), .B1(n31589), .Y(
        n18455) );
  AOI22XL U22941 ( .A0(n16666), .A1(conv_3[380]), .B0(n16662), .B1(conv_3[395]), .Y(n18458) );
  NAND2XL U22942 ( .A(n18458), .B(n18457), .Y(n26191) );
  INVXL U22943 ( .A(conv_3[185]), .Y(n31619) );
  INVXL U22944 ( .A(conv_3[215]), .Y(n28830) );
  INVXL U22945 ( .A(conv_3[230]), .Y(n29160) );
  OAI22XL U22946 ( .A0(n22612), .A1(n28830), .B0(n18321), .B1(n29160), .Y(
        n18459) );
  AOI211XL U22947 ( .A0(conv_3[200]), .A1(n22762), .B0(n18460), .C0(n18459), 
        .Y(n28310) );
  INVXL U22948 ( .A(n28310), .Y(n35046) );
  AOI22XL U22949 ( .A0(n16667), .A1(n26191), .B0(n16670), .B1(n35046), .Y(
        n18467) );
  AOI22XL U22950 ( .A0(n25306), .A1(conv_3[320]), .B0(n16662), .B1(conv_3[335]), .Y(n18462) );
  AOI22XL U22951 ( .A0(n18658), .A1(conv_3[305]), .B0(n16673), .B1(conv_3[350]), .Y(n18461) );
  NAND2XL U22952 ( .A(n18462), .B(n18461), .Y(n26192) );
  AOI22XL U22953 ( .A0(n16662), .A1(conv_3[95]), .B0(n22690), .B1(conv_3[65]), 
        .Y(n18464) );
  NAND2XL U22954 ( .A(n18465), .B(n18464), .Y(n35052) );
  AOI22XL U22955 ( .A0(n16659), .A1(n26192), .B0(n18463), .B1(n35052), .Y(
        n18466) );
  OAI211XL U22956 ( .A0(n35041), .A1(n26621), .B0(n18467), .C0(n18466), .Y(
        n18468) );
  NOR3XL U22957 ( .A(n18470), .B(n18469), .C(n18468), .Y(n18708) );
  AOI22XL U22958 ( .A0(n16666), .A1(conv_3[383]), .B0(n16673), .B1(conv_3[413]), .Y(n18472) );
  AOI22XL U22959 ( .A0(n16662), .A1(conv_3[398]), .B0(n22616), .B1(conv_3[368]), .Y(n18471) );
  NAND2XL U22960 ( .A(n18472), .B(n18471), .Y(n26244) );
  INVXL U22961 ( .A(conv_3[263]), .Y(n32100) );
  INVXL U22962 ( .A(conv_3[248]), .Y(n35695) );
  AOI22XL U22963 ( .A0(n20735), .A1(n32100), .B0(n35695), .B1(n18634), .Y(
        n21333) );
  AOI222XL U22964 ( .A0(n21333), .A1(n22713), .B0(n16673), .B1(conv_3[293]), 
        .C0(conv_3[278]), .C1(n25289), .Y(n35030) );
  INVXL U22965 ( .A(conv_3[188]), .Y(n31595) );
  INVXL U22966 ( .A(conv_3[218]), .Y(n32061) );
  INVXL U22967 ( .A(conv_3[233]), .Y(n35675) );
  OAI22XL U22968 ( .A0(n22612), .A1(n32061), .B0(n24039), .B1(n35675), .Y(
        n18473) );
  AOI211XL U22969 ( .A0(conv_3[203]), .A1(n22762), .B0(n18474), .C0(n18473), 
        .Y(n35033) );
  INVX2 U22970 ( .A(n18475), .Y(n28553) );
  OAI22XL U22971 ( .A0(n35030), .A1(n28575), .B0(n35033), .B1(n28553), .Y(
        n18488) );
  INVXL U22972 ( .A(conv_3[473]), .Y(n33014) );
  INVXL U22973 ( .A(conv_3[458]), .Y(n35804) );
  AOI22XL U22974 ( .A0(n20735), .A1(n33014), .B0(n35804), .B1(n19855), .Y(
        n21340) );
  AOI222XL U22975 ( .A0(n21340), .A1(n36246), .B0(n22759), .B1(conv_3[428]), 
        .C0(n16666), .C1(conv_3[443]), .Y(n25732) );
  INVXL U22976 ( .A(n25732), .Y(n35031) );
  AOI22XL U22977 ( .A0(n20735), .A1(conv_3[533]), .B0(conv_3[518]), .B1(n18526), .Y(n20513) );
  AOI22XL U22978 ( .A0(n20735), .A1(conv_3[503]), .B0(conv_3[488]), .B1(n18516), .Y(n20514) );
  AOI22XL U22979 ( .A0(n26263), .A1(n35031), .B0(n28571), .B1(n35034), .Y(
        n18486) );
  INVXL U22980 ( .A(conv_3[53]), .Y(n34393) );
  INVXL U22981 ( .A(conv_3[23]), .Y(n31272) );
  INVXL U22982 ( .A(conv_3[38]), .Y(n35593) );
  OAI22XL U22983 ( .A0(n19902), .A1(n31272), .B0(n22612), .B1(n35593), .Y(
        n18476) );
  AOI211XL U22984 ( .A0(conv_3[8]), .A1(n22759), .B0(n18477), .C0(n18476), .Y(
        n26246) );
  INVXL U22985 ( .A(n26246), .Y(n35032) );
  AOI22XL U22986 ( .A0(n25306), .A1(conv_3[143]), .B0(n16673), .B1(conv_3[173]), .Y(n18479) );
  AOI22XL U22987 ( .A0(n16662), .A1(conv_3[158]), .B0(n22759), .B1(conv_3[128]), .Y(n18478) );
  NAND2XL U22988 ( .A(n18479), .B(n18478), .Y(n28344) );
  AOI22XL U22989 ( .A0(n16660), .A1(n35032), .B0(n28324), .B1(n28344), .Y(
        n18485) );
  AOI22XL U22990 ( .A0(n16662), .A1(conv_3[338]), .B0(n22616), .B1(conv_3[308]), .Y(n18481) );
  AOI22XL U22991 ( .A0(n16666), .A1(conv_3[323]), .B0(n16673), .B1(conv_3[353]), .Y(n18480) );
  NAND2XL U22992 ( .A(n18481), .B(n18480), .Y(n26245) );
  AOI22XL U22993 ( .A0(n16666), .A1(conv_3[83]), .B0(n16673), .B1(conv_3[113]), 
        .Y(n18483) );
  AOI22XL U22994 ( .A0(n16662), .A1(conv_3[98]), .B0(n22616), .B1(conv_3[68]), 
        .Y(n18482) );
  NAND2XL U22995 ( .A(n18483), .B(n18482), .Y(n35040) );
  AOI22XL U22996 ( .A0(n16659), .A1(n26245), .B0(n18463), .B1(n35040), .Y(
        n18484) );
  NAND3XL U22997 ( .A(n18486), .B(n18485), .C(n18484), .Y(n18487) );
  AOI211XL U22998 ( .A0(n16667), .A1(n26244), .B0(n18488), .C0(n18487), .Y(
        n18707) );
  AOI22XL U22999 ( .A0(n22762), .A1(conv_3[139]), .B0(n16662), .B1(conv_3[154]), .Y(n18489) );
  NAND2XL U23000 ( .A(n18490), .B(n18489), .Y(n35102) );
  AOI22XL U23001 ( .A0(n20735), .A1(conv_3[529]), .B0(conv_3[514]), .B1(n19253), .Y(n20495) );
  AOI22XL U23002 ( .A0(n20735), .A1(conv_3[499]), .B0(conv_3[484]), .B1(n19253), .Y(n20490) );
  INVXL U23003 ( .A(n22770), .Y(n18776) );
  INVXL U23004 ( .A(conv_3[199]), .Y(n22150) );
  INVXL U23005 ( .A(conv_3[214]), .Y(n23627) );
  INVXL U23006 ( .A(conv_3[229]), .Y(n22168) );
  OAI22XL U23007 ( .A0(n22612), .A1(n23627), .B0(n24039), .B1(n22168), .Y(
        n18491) );
  AOI211XL U23008 ( .A0(conv_3[184]), .A1(n22759), .B0(n18492), .C0(n18491), 
        .Y(n24827) );
  AOI211XL U23009 ( .A0(n28407), .A1(n35102), .B0(n18498), .C0(n18493), .Y(
        n25763) );
  AOI22XL U23010 ( .A0(n22762), .A1(conv_3[19]), .B0(n16662), .B1(conv_3[34]), 
        .Y(n18494) );
  NAND2XL U23011 ( .A(n18495), .B(n18494), .Y(n26208) );
  INVXL U23012 ( .A(conv_3[94]), .Y(n22881) );
  INVXL U23013 ( .A(conv_3[64]), .Y(n23904) );
  INVXL U23014 ( .A(conv_3[109]), .Y(n22915) );
  OAI22XL U23015 ( .A0(n22550), .A1(n23904), .B0(n24039), .B1(n22915), .Y(
        n18496) );
  AOI211XL U23016 ( .A0(conv_3[79]), .A1(n22762), .B0(n18497), .C0(n18496), 
        .Y(n35107) );
  AOI211XL U23017 ( .A0(n21100), .A1(n26208), .B0(n18499), .C0(n18498), .Y(
        n25762) );
  INVXL U23018 ( .A(conv_3[469]), .Y(n22195) );
  INVXL U23019 ( .A(conv_3[454]), .Y(n24265) );
  AOI22XL U23020 ( .A0(n20735), .A1(n22195), .B0(n24265), .B1(n18634), .Y(
        n21201) );
  AOI222XL U23021 ( .A0(n21201), .A1(n36246), .B0(n22690), .B1(conv_3[424]), 
        .C0(n22762), .C1(conv_3[439]), .Y(n25770) );
  NAND2XL U23022 ( .A(N18014), .B(n22369), .Y(n25393) );
  AOI22XL U23023 ( .A0(n22762), .A1(conv_3[379]), .B0(n16662), .B1(conv_3[394]), .Y(n18500) );
  NAND2XL U23024 ( .A(n18501), .B(n18500), .Y(n25767) );
  OAI2BB2XL U23025 ( .B0(n25770), .B1(n25393), .A0N(n25399), .A1N(n25767), .Y(
        n18505) );
  INVXL U23026 ( .A(conv_3[304]), .Y(n23227) );
  INVXL U23027 ( .A(conv_3[319]), .Y(n23815) );
  INVXL U23028 ( .A(conv_3[334]), .Y(n26950) );
  OAI22XL U23029 ( .A0(n19902), .A1(n23815), .B0(n22612), .B1(n26950), .Y(
        n18502) );
  AOI211XL U23030 ( .A0(conv_3[349]), .A1(n16723), .B0(n18503), .C0(n18502), 
        .Y(n25761) );
  INVXL U23031 ( .A(n28289), .Y(n25395) );
  INVXL U23032 ( .A(conv_3[259]), .Y(n22117) );
  INVXL U23033 ( .A(conv_3[244]), .Y(n24030) );
  AOI22XL U23034 ( .A0(n20735), .A1(n22117), .B0(n24030), .B1(n18526), .Y(
        n21195) );
  AOI222XL U23035 ( .A0(n21195), .A1(n22713), .B0(n16673), .B1(conv_3[289]), 
        .C0(conv_3[274]), .C1(n25289), .Y(n35103) );
  NOR2XL U23036 ( .A(N18014), .B(n19181), .Y(n25337) );
  OAI22XL U23037 ( .A0(n25761), .A1(n25395), .B0(n35103), .B1(n25402), .Y(
        n18504) );
  AOI211XL U23038 ( .A0(n36244), .A1(n35104), .B0(n18505), .C0(n18504), .Y(
        n26210) );
  OAI222XL U23039 ( .A0(n35135), .A1(n25763), .B0(n34989), .B1(n25762), .C0(
        n26210), .C1(N18471), .Y(n18723) );
  AOI22XL U23040 ( .A0(n20735), .A1(conv_3[475]), .B0(conv_3[460]), .B1(n18526), .Y(n19436) );
  INVXL U23041 ( .A(n19436), .Y(n21353) );
  AOI222XL U23042 ( .A0(conv_3[430]), .A1(n22759), .B0(n36246), .B1(n21353), 
        .C0(n22762), .C1(conv_3[445]), .Y(n35056) );
  INVXL U23043 ( .A(n35056), .Y(n28352) );
  AOI22XL U23044 ( .A0(n16666), .A1(conv_3[145]), .B0(n18240), .B1(conv_3[175]), .Y(n18507) );
  AOI22XL U23045 ( .A0(n16662), .A1(conv_3[160]), .B0(n22759), .B1(conv_3[130]), .Y(n18506) );
  NAND2XL U23046 ( .A(n18507), .B(n18506), .Y(n28351) );
  AOI22XL U23047 ( .A0(n26263), .A1(n28352), .B0(n28324), .B1(n28351), .Y(
        n18523) );
  AOI22XL U23048 ( .A0(n25299), .A1(conv_3[310]), .B0(n18240), .B1(conv_3[355]), .Y(n18509) );
  NAND2XL U23049 ( .A(n18509), .B(n18508), .Y(n26240) );
  AOI22XL U23050 ( .A0(n16666), .A1(conv_3[385]), .B0(n16673), .B1(conv_3[415]), .Y(n18511) );
  AOI22XL U23051 ( .A0(n16662), .A1(conv_3[400]), .B0(n22759), .B1(conv_3[370]), .Y(n18510) );
  NAND2XL U23052 ( .A(n18511), .B(n18510), .Y(n26237) );
  AOI22XL U23053 ( .A0(n28528), .A1(n26240), .B0(n16667), .B1(n26237), .Y(
        n18522) );
  AOI22XL U23054 ( .A0(n20735), .A1(conv_3[535]), .B0(conv_3[520]), .B1(n19253), .Y(n21357) );
  AOI22XL U23055 ( .A0(n20735), .A1(conv_3[505]), .B0(conv_3[490]), .B1(n18516), .Y(n21359) );
  INVXL U23056 ( .A(conv_3[70]), .Y(n31435) );
  INVXL U23057 ( .A(conv_3[85]), .Y(n31809) );
  INVXL U23058 ( .A(conv_3[100]), .Y(n31672) );
  OAI22XL U23059 ( .A0(n19902), .A1(n31809), .B0(n22612), .B1(n31672), .Y(
        n18512) );
  AOI211XL U23060 ( .A0(n16673), .A1(conv_3[115]), .B0(n18513), .C0(n18512), 
        .Y(n25726) );
  INVXL U23061 ( .A(conv_3[40]), .Y(n31237) );
  INVXL U23062 ( .A(conv_3[25]), .Y(n31256) );
  INVXL U23063 ( .A(conv_3[55]), .Y(n31203) );
  OAI22XL U23064 ( .A0(n22546), .A1(n31256), .B0(n18321), .B1(n31203), .Y(
        n18514) );
  OAI22XL U23065 ( .A0(n25726), .A1(n16672), .B0(n35055), .B1(n35198), .Y(
        n18520) );
  OAI22XL U23066 ( .A0(n18516), .A1(conv_3[265]), .B0(conv_3[250]), .B1(n35269), .Y(n19427) );
  AOI222XL U23067 ( .A0(n21371), .A1(n22765), .B0(n16673), .B1(conv_3[295]), 
        .C0(conv_3[280]), .C1(n16662), .Y(n35053) );
  INVXL U23068 ( .A(conv_3[235]), .Y(n29166) );
  INVXL U23069 ( .A(conv_3[220]), .Y(n31535) );
  INVXL U23070 ( .A(conv_3[190]), .Y(n31613) );
  OAI22XL U23071 ( .A0(n22612), .A1(n31535), .B0(n16668), .B1(n31613), .Y(
        n18517) );
  AOI211XL U23072 ( .A0(conv_3[205]), .A1(n22762), .B0(n18518), .C0(n18517), 
        .Y(n35057) );
  OAI22XL U23073 ( .A0(n35053), .A1(n28575), .B0(n35057), .B1(n28553), .Y(
        n18519) );
  AOI211XL U23074 ( .A0(n28571), .A1(n35054), .B0(n18520), .C0(n18519), .Y(
        n18521) );
  NAND3XL U23075 ( .A(n18523), .B(n18522), .C(n18521), .Y(n18712) );
  AOI22XL U23076 ( .A0(n16666), .A1(conv_3[22]), .B0(n22759), .B1(conv_3[7]), 
        .Y(n18525) );
  NAND2XL U23077 ( .A(n18525), .B(n18524), .Y(n35094) );
  INVXL U23078 ( .A(conv_3[532]), .Y(n27571) );
  INVXL U23079 ( .A(conv_3[517]), .Y(n31166) );
  AOI22XL U23080 ( .A0(n20735), .A1(n27571), .B0(n31166), .B1(n18634), .Y(
        n21226) );
  INVXL U23081 ( .A(conv_3[502]), .Y(n32064) );
  INVXL U23082 ( .A(conv_3[487]), .Y(n35825) );
  AOI22XL U23083 ( .A0(n35269), .A1(n32064), .B0(n35825), .B1(n18526), .Y(
        n21213) );
  INVXL U23084 ( .A(conv_3[262]), .Y(n29111) );
  INVXL U23085 ( .A(conv_3[247]), .Y(n35688) );
  AOI22XL U23086 ( .A0(n20735), .A1(n29111), .B0(n35688), .B1(n18526), .Y(
        n21228) );
  AOI222XL U23087 ( .A0(n21228), .A1(n22743), .B0(n16673), .B1(conv_3[292]), 
        .C0(conv_3[277]), .C1(n25289), .Y(n28315) );
  OAI22XL U23088 ( .A0(n28551), .A1(n35090), .B0(n28315), .B1(n34981), .Y(
        n18542) );
  INVXL U23089 ( .A(conv_3[472]), .Y(n32338) );
  INVXL U23090 ( .A(conv_3[457]), .Y(n33782) );
  AOI22XL U23091 ( .A0(n20735), .A1(n32338), .B0(n33782), .B1(n18526), .Y(
        n21217) );
  AOI222XL U23092 ( .A0(n21217), .A1(n36246), .B0(n22759), .B1(conv_3[427]), 
        .C0(n25306), .C1(conv_3[442]), .Y(n35089) );
  AOI22XL U23093 ( .A0(n16662), .A1(conv_3[397]), .B0(n22759), .B1(conv_3[367]), .Y(n18527) );
  NAND2XL U23094 ( .A(n18528), .B(n18527), .Y(n26214) );
  AOI22XL U23095 ( .A0(n26263), .A1(n26216), .B0(n16667), .B1(n26214), .Y(
        n18540) );
  AOI22XL U23096 ( .A0(n16666), .A1(conv_3[202]), .B0(n22759), .B1(conv_3[187]), .Y(n18529) );
  NAND2XL U23097 ( .A(n18530), .B(n18529), .Y(n35100) );
  INVXL U23098 ( .A(conv_3[97]), .Y(n31678) );
  INVXL U23099 ( .A(conv_3[82]), .Y(n31838) );
  INVXL U23100 ( .A(conv_3[112]), .Y(n31802) );
  OAI22XL U23101 ( .A0(n19401), .A1(n31838), .B0(n18321), .B1(n31802), .Y(
        n18531) );
  AOI211XL U23102 ( .A0(conv_3[67]), .A1(n22759), .B0(n18532), .C0(n18531), 
        .Y(n26213) );
  INVXL U23103 ( .A(n26213), .Y(n35092) );
  AOI22XL U23104 ( .A0(n16665), .A1(n35100), .B0(n18463), .B1(n35092), .Y(
        n18539) );
  AOI22XL U23105 ( .A0(n18658), .A1(conv_3[307]), .B0(n16673), .B1(conv_3[352]), .Y(n18534) );
  AOI22XL U23106 ( .A0(n16666), .A1(conv_3[322]), .B0(n16662), .B1(conv_3[337]), .Y(n18533) );
  NAND2XL U23107 ( .A(n18534), .B(n18533), .Y(n26215) );
  AOI22XL U23108 ( .A0(n16662), .A1(conv_3[157]), .B0(n22759), .B1(conv_3[127]), .Y(n18536) );
  NAND2XL U23109 ( .A(n18537), .B(n18536), .Y(n35091) );
  AOI22XL U23110 ( .A0(n28528), .A1(n26215), .B0(n28324), .B1(n35091), .Y(
        n18538) );
  NAND3XL U23111 ( .A(n18540), .B(n18539), .C(n18538), .Y(n18541) );
  AOI211XL U23112 ( .A0(n16660), .A1(n35094), .B0(n18542), .C0(n18541), .Y(
        n18706) );
  AOI22XL U23113 ( .A0(n16666), .A1(conv_3[381]), .B0(n16662), .B1(conv_3[396]), .Y(n18543) );
  NAND2XL U23114 ( .A(n18544), .B(n18543), .Y(n26200) );
  INVXL U23115 ( .A(conv_3[531]), .Y(n26307) );
  INVXL U23116 ( .A(conv_3[516]), .Y(n31177) );
  AOI22XL U23117 ( .A0(n20735), .A1(n26307), .B0(n31177), .B1(n19253), .Y(
        n21263) );
  INVXL U23118 ( .A(conv_3[501]), .Y(n35840) );
  AOI2BB2XL U23119 ( .B0(n20735), .B1(n35840), .A0N(conv_3[486]), .A1N(n35269), 
        .Y(n21269) );
  INVXL U23120 ( .A(conv_3[261]), .Y(n29135) );
  INVXL U23121 ( .A(conv_3[246]), .Y(n35682) );
  AOI22XL U23122 ( .A0(n20735), .A1(n29135), .B0(n35682), .B1(n18526), .Y(
        n21265) );
  AOI222XL U23123 ( .A0(n21265), .A1(n22743), .B0(n16673), .B1(conv_3[291]), 
        .C0(conv_3[276]), .C1(n25289), .Y(n35065) );
  AOI22XL U23124 ( .A0(n25306), .A1(conv_3[201]), .B0(n18240), .B1(conv_3[231]), .Y(n18546) );
  AOI22XL U23125 ( .A0(n16662), .A1(conv_3[216]), .B0(n22690), .B1(conv_3[186]), .Y(n18545) );
  NAND2XL U23126 ( .A(n18546), .B(n18545), .Y(n35069) );
  AOI22XL U23127 ( .A0(n25306), .A1(conv_3[81]), .B0(n22759), .B1(conv_3[66]), 
        .Y(n18547) );
  NAND2XL U23128 ( .A(n18548), .B(n18547), .Y(n35073) );
  AOI22XL U23129 ( .A0(n16665), .A1(n35069), .B0(n18463), .B1(n35073), .Y(
        n18558) );
  AOI22XL U23130 ( .A0(n16662), .A1(conv_3[336]), .B0(n22759), .B1(conv_3[306]), .Y(n18549) );
  NAND2XL U23131 ( .A(n18550), .B(n18549), .Y(n26199) );
  INVXL U23132 ( .A(conv_3[36]), .Y(n31249) );
  INVXL U23133 ( .A(conv_3[21]), .Y(n31278) );
  INVXL U23134 ( .A(conv_3[51]), .Y(n31215) );
  OAI22XL U23135 ( .A0(n22546), .A1(n31278), .B0(n24039), .B1(n31215), .Y(
        n18551) );
  AOI211XL U23136 ( .A0(conv_3[6]), .A1(n22616), .B0(n18552), .C0(n18551), .Y(
        n35068) );
  INVXL U23137 ( .A(conv_3[471]), .Y(n35812) );
  INVXL U23138 ( .A(conv_3[456]), .Y(n31512) );
  AOI22XL U23139 ( .A0(n20735), .A1(n35812), .B0(n31512), .B1(n18634), .Y(
        n21270) );
  AOI222XL U23140 ( .A0(n21270), .A1(n36246), .B0(n22759), .B1(conv_3[426]), 
        .C0(n25306), .C1(conv_3[441]), .Y(n28321) );
  INVXL U23141 ( .A(conv_3[141]), .Y(n31718) );
  INVXL U23142 ( .A(conv_3[156]), .Y(n32313) );
  INVXL U23143 ( .A(conv_3[171]), .Y(n31566) );
  OAI22XL U23144 ( .A0(n22612), .A1(n32313), .B0(n24039), .B1(n31566), .Y(
        n18553) );
  AOI211XL U23145 ( .A0(conv_3[126]), .A1(n22616), .B0(n18554), .C0(n18553), 
        .Y(n35067) );
  OAI22XL U23146 ( .A0(n28321), .A1(n34958), .B0(n35067), .B1(n26621), .Y(
        n18555) );
  AOI211XL U23147 ( .A0(n34992), .A1(n26199), .B0(n18556), .C0(n18555), .Y(
        n18557) );
  OAI211XL U23148 ( .A0(n35065), .A1(n28575), .B0(n18558), .C0(n18557), .Y(
        n18559) );
  AOI211XL U23149 ( .A0(n16667), .A1(n26200), .B0(n18560), .C0(n18559), .Y(
        n18717) );
  AOI22XL U23150 ( .A0(n25299), .A1(conv_3[69]), .B0(n16673), .B1(conv_3[114]), 
        .Y(n18562) );
  AOI22XL U23151 ( .A0(n20978), .A1(conv_3[84]), .B0(n16662), .B1(conv_3[99]), 
        .Y(n18561) );
  NAND2XL U23152 ( .A(n18562), .B(n18561), .Y(n35082) );
  INVXL U23153 ( .A(n35082), .Y(n28332) );
  INVXL U23154 ( .A(conv_3[399]), .Y(n32047) );
  INVXL U23155 ( .A(conv_3[414]), .Y(n32555) );
  OAI22XL U23156 ( .A0(n22612), .A1(n32047), .B0(n18321), .B1(n32555), .Y(
        n18564) );
  INVXL U23157 ( .A(conv_3[384]), .Y(n31506) );
  INVXL U23158 ( .A(conv_3[369]), .Y(n35763) );
  OAI22XL U23159 ( .A0(n19902), .A1(n31506), .B0(n22717), .B1(n35763), .Y(
        n18563) );
  OAI22XL U23160 ( .A0(n28332), .A1(n16672), .B0(n26223), .B1(n28577), .Y(
        n18577) );
  INVXL U23161 ( .A(conv_3[219]), .Y(n31541) );
  INVXL U23162 ( .A(conv_3[234]), .Y(n30694) );
  OAI22XL U23163 ( .A0(n22612), .A1(n31541), .B0(n18321), .B1(n30694), .Y(
        n18566) );
  INVXL U23164 ( .A(conv_3[204]), .Y(n31847) );
  INVXL U23165 ( .A(conv_3[189]), .Y(n31608) );
  OAI22XL U23166 ( .A0(n19902), .A1(n31847), .B0(n22717), .B1(n31608), .Y(
        n18565) );
  AOI22XL U23167 ( .A0(n16662), .A1(conv_3[339]), .B0(n22616), .B1(conv_3[309]), .Y(n18568) );
  NAND2XL U23168 ( .A(n18568), .B(n18567), .Y(n26222) );
  INVXL U23169 ( .A(n26222), .Y(n24864) );
  OAI22XL U23170 ( .A0(n35085), .A1(n28553), .B0(n24864), .B1(n28479), .Y(
        n18576) );
  INVXL U23171 ( .A(conv_3[534]), .Y(n28961) );
  INVXL U23172 ( .A(conv_3[519]), .Y(n31152) );
  AOI22XL U23173 ( .A0(n20735), .A1(n28961), .B0(n31152), .B1(n18526), .Y(
        n21295) );
  INVXL U23174 ( .A(conv_3[504]), .Y(n32081) );
  INVXL U23175 ( .A(conv_3[489]), .Y(n31549) );
  AOI22XL U23176 ( .A0(n20735), .A1(n32081), .B0(n31549), .B1(n18526), .Y(
        n21286) );
  INVXL U23177 ( .A(conv_3[474]), .Y(n33018) );
  AOI2BB2XL U23178 ( .B0(n20735), .B1(n33018), .A0N(conv_3[459]), .A1N(n35269), 
        .Y(n21282) );
  AOI222XL U23179 ( .A0(n21282), .A1(n36246), .B0(n22759), .B1(conv_3[429]), 
        .C0(n25306), .C1(conv_3[444]), .Y(n35078) );
  INVXL U23180 ( .A(n35078), .Y(n28330) );
  AOI22XL U23181 ( .A0(n22759), .A1(conv_3[129]), .B0(n18240), .B1(conv_3[174]), .Y(n18569) );
  NAND2XL U23182 ( .A(n18570), .B(n18569), .Y(n35079) );
  AOI22XL U23183 ( .A0(n26263), .A1(n28330), .B0(n28366), .B1(n35079), .Y(
        n18574) );
  INVXL U23184 ( .A(conv_3[264]), .Y(n32106) );
  INVXL U23185 ( .A(conv_3[249]), .Y(n35702) );
  AOI22XL U23186 ( .A0(n20735), .A1(n32106), .B0(n35702), .B1(n18516), .Y(
        n21297) );
  AOI222XL U23187 ( .A0(n21297), .A1(n22713), .B0(n18810), .B1(conv_3[279]), 
        .C0(conv_3[294]), .C1(n16673), .Y(n35077) );
  INVXL U23188 ( .A(n35077), .Y(n28329) );
  AOI22XL U23189 ( .A0(n20978), .A1(conv_3[24]), .B0(n18240), .B1(conv_3[54]), 
        .Y(n18572) );
  AOI22XL U23190 ( .A0(n16662), .A1(conv_3[39]), .B0(n22616), .B1(conv_3[9]), 
        .Y(n18571) );
  NAND2XL U23191 ( .A(n18572), .B(n18571), .Y(n35080) );
  AOI22XL U23192 ( .A0(n28414), .A1(n28329), .B0(n18197), .B1(n35080), .Y(
        n18573) );
  OAI211XL U23193 ( .A0(n28551), .A1(n35081), .B0(n18574), .C0(n18573), .Y(
        n18575) );
  NOR3XL U23194 ( .A(n18577), .B(n18576), .C(n18575), .Y(n18716) );
  AOI22XL U23195 ( .A0(n20735), .A1(conv_3[536]), .B0(conv_3[521]), .B1(n19253), .Y(n21313) );
  AOI22XL U23196 ( .A0(n20735), .A1(conv_3[506]), .B0(conv_3[491]), .B1(n18634), .Y(n20473) );
  INVXL U23197 ( .A(n35114), .Y(n24859) );
  AOI22XL U23198 ( .A0(n16662), .A1(conv_3[221]), .B0(n22759), .B1(conv_3[191]), .Y(n18579) );
  AOI22XL U23199 ( .A0(n16666), .A1(conv_3[206]), .B0(n18240), .B1(conv_3[236]), .Y(n18578) );
  NAND2XL U23200 ( .A(n18579), .B(n18578), .Y(n25754) );
  INVXL U23201 ( .A(n25754), .Y(n35113) );
  OAI22XL U23202 ( .A0(n28551), .A1(n24859), .B0(n35113), .B1(n28553), .Y(
        n18594) );
  INVXL U23203 ( .A(conv_3[131]), .Y(n31442) );
  INVXL U23204 ( .A(conv_3[146]), .Y(n33971) );
  INVXL U23205 ( .A(conv_3[161]), .Y(n32320) );
  OAI22XL U23206 ( .A0(n19401), .A1(n33971), .B0(n22612), .B1(n32320), .Y(
        n18580) );
  AOI211XL U23207 ( .A0(conv_3[176]), .A1(n16673), .B0(n18581), .C0(n18580), 
        .Y(n28339) );
  INVXL U23208 ( .A(conv_3[476]), .Y(n32344) );
  INVXL U23209 ( .A(conv_3[461]), .Y(n31528) );
  AOI22XL U23210 ( .A0(n20735), .A1(n32344), .B0(n31528), .B1(n18526), .Y(
        n21314) );
  AOI222XL U23211 ( .A0(n21314), .A1(n36246), .B0(n22759), .B1(conv_3[431]), 
        .C0(n22762), .C1(conv_3[446]), .Y(n35112) );
  OAI22XL U23212 ( .A0(n28339), .A1(n26621), .B0(n35112), .B1(n34958), .Y(
        n18593) );
  INVXL U23213 ( .A(conv_3[416]), .Y(n32015) );
  INVXL U23214 ( .A(conv_3[401]), .Y(n32042) );
  INVXL U23215 ( .A(conv_3[371]), .Y(n31635) );
  OAI22XL U23216 ( .A0(n22612), .A1(n32042), .B0(n22717), .B1(n31635), .Y(
        n18582) );
  AOI211XL U23217 ( .A0(conv_3[386]), .A1(n16666), .B0(n18583), .C0(n18582), 
        .Y(n26229) );
  AOI22XL U23218 ( .A0(n16662), .A1(conv_3[41]), .B0(n22759), .B1(conv_3[11]), 
        .Y(n18585) );
  AOI22XL U23219 ( .A0(n16666), .A1(conv_3[26]), .B0(n16673), .B1(conv_3[56]), 
        .Y(n18584) );
  NAND2XL U23220 ( .A(n18585), .B(n18584), .Y(n35123) );
  AOI22XL U23221 ( .A0(n22759), .A1(conv_3[71]), .B0(n16673), .B1(conv_3[116]), 
        .Y(n18587) );
  AOI22XL U23222 ( .A0(n16666), .A1(conv_3[86]), .B0(n16662), .B1(conv_3[101]), 
        .Y(n18586) );
  NAND2XL U23223 ( .A(n18587), .B(n18586), .Y(n35115) );
  AOI22XL U23224 ( .A0(n16660), .A1(n35123), .B0(n18463), .B1(n35115), .Y(
        n18591) );
  AOI22XL U23225 ( .A0(n16666), .A1(conv_3[326]), .B0(n16673), .B1(conv_3[356]), .Y(n18589) );
  AOI22XL U23226 ( .A0(n16662), .A1(conv_3[341]), .B0(n22616), .B1(conv_3[311]), .Y(n18588) );
  NAND2XL U23227 ( .A(n18589), .B(n18588), .Y(n26232) );
  OAI22XL U23228 ( .A0(n18526), .A1(conv_3[266]), .B0(conv_3[251]), .B1(n35269), .Y(n21312) );
  INVXL U23229 ( .A(n21312), .Y(n21318) );
  AOI222XL U23230 ( .A0(n21318), .A1(n22743), .B0(n16673), .B1(conv_3[296]), 
        .C0(conv_3[281]), .C1(n25289), .Y(n25755) );
  INVXL U23231 ( .A(n25755), .Y(n35116) );
  OAI211XL U23232 ( .A0(n26229), .A1(n28577), .B0(n18591), .C0(n18590), .Y(
        n18592) );
  NOR3XL U23233 ( .A(n18594), .B(n18593), .C(n18592), .Y(n18711) );
  NAND4XL U23234 ( .A(n18706), .B(n18717), .C(n18716), .D(n18711), .Y(n18595)
         );
  NOR3XL U23235 ( .A(n18723), .B(n18712), .C(n18595), .Y(n18596) );
  AOI31XL U23236 ( .A0(n18708), .A1(n18707), .A2(n18596), .B0(pool[119]), .Y(
        n18653) );
  AOI22XL U23237 ( .A0(n20735), .A1(conv_3[528]), .B0(conv_3[513]), .B1(n19253), .Y(n20422) );
  AOI22XL U23238 ( .A0(n20735), .A1(conv_3[498]), .B0(conv_3[483]), .B1(n18634), .Y(n21123) );
  INVXL U23239 ( .A(n26171), .Y(n35133) );
  AOI22XL U23240 ( .A0(n18658), .A1(conv_3[183]), .B0(n18240), .B1(conv_3[228]), .Y(n18597) );
  NAND2XL U23241 ( .A(n18598), .B(n18597), .Y(n35128) );
  AOI22XL U23242 ( .A0(n25306), .A1(conv_3[138]), .B0(n16662), .B1(conv_3[153]), .Y(n18599) );
  NAND2XL U23243 ( .A(n18600), .B(n18599), .Y(n35127) );
  AOI22XL U23244 ( .A0(n22362), .A1(n35128), .B0(n28407), .B1(n35127), .Y(
        n18601) );
  NAND2BXL U23245 ( .AN(n25701), .B(n18601), .Y(n25706) );
  AOI22XL U23246 ( .A0(n25306), .A1(conv_3[378]), .B0(n16662), .B1(conv_3[393]), .Y(n18603) );
  AOI22XL U23247 ( .A0(n18658), .A1(conv_3[363]), .B0(n18240), .B1(conv_3[408]), .Y(n18602) );
  NAND2XL U23248 ( .A(n18603), .B(n18602), .Y(n25699) );
  AOI22XL U23249 ( .A0(n25306), .A1(conv_3[318]), .B0(n22759), .B1(conv_3[303]), .Y(n18605) );
  AOI22XL U23250 ( .A0(n16662), .A1(conv_3[333]), .B0(n16723), .B1(conv_3[348]), .Y(n18604) );
  NAND2XL U23251 ( .A(n18605), .B(n18604), .Y(n25700) );
  NAND2XL U23252 ( .A(n36244), .B(n26171), .Y(n24848) );
  OAI2BB1XL U23253 ( .A0N(n28289), .A1N(n25700), .B0(n24848), .Y(n18607) );
  INVXL U23254 ( .A(conv_3[258]), .Y(n29419) );
  INVXL U23255 ( .A(conv_3[243]), .Y(n29662) );
  AOI22XL U23256 ( .A0(n20735), .A1(n29419), .B0(n29662), .B1(n19253), .Y(
        n21130) );
  AOI222XL U23257 ( .A0(n21130), .A1(n22743), .B0(n16673), .B1(conv_3[288]), 
        .C0(conv_3[273]), .C1(n25289), .Y(n25698) );
  INVXL U23258 ( .A(conv_3[468]), .Y(n30189) );
  AOI222XL U23259 ( .A0(n21124), .A1(n36246), .B0(n22690), .B1(conv_3[423]), 
        .C0(n22770), .C1(conv_3[438]), .Y(n25697) );
  OAI22XL U23260 ( .A0(n25698), .A1(n25402), .B0(n25697), .B1(n25393), .Y(
        n18606) );
  AOI22XL U23261 ( .A0(n16662), .A1(conv_3[33]), .B0(n16673), .B1(conv_3[48]), 
        .Y(n18609) );
  AOI22XL U23262 ( .A0(n25306), .A1(conv_3[18]), .B0(n25299), .B1(conv_3[3]), 
        .Y(n18608) );
  NAND2XL U23263 ( .A(n18609), .B(n18608), .Y(n26170) );
  INVXL U23264 ( .A(conv_3[108]), .Y(n29655) );
  INVXL U23265 ( .A(conv_3[93]), .Y(n29642) );
  INVXL U23266 ( .A(conv_3[63]), .Y(n34112) );
  OAI22XL U23267 ( .A0(n22612), .A1(n29642), .B0(n22717), .B1(n34112), .Y(
        n18610) );
  AOI211XL U23268 ( .A0(n21100), .A1(n26170), .B0(n18612), .C0(n25701), .Y(
        n25703) );
  OAI22XL U23269 ( .A0(N18471), .A1(n26175), .B0(n25703), .B1(n34989), .Y(
        n18613) );
  INVXL U23270 ( .A(pool[117]), .Y(n24568) );
  AOI22XL U23271 ( .A0(n20735), .A1(conv_3[527]), .B0(conv_3[512]), .B1(n18526), .Y(n19470) );
  AOI22XL U23272 ( .A0(n20735), .A1(conv_3[497]), .B0(conv_3[482]), .B1(n19253), .Y(n20432) );
  INVXL U23273 ( .A(n28278), .Y(n35142) );
  AOI22XL U23274 ( .A0(n20735), .A1(conv_3[257]), .B0(conv_3[242]), .B1(n18526), .Y(n19471) );
  INVXL U23275 ( .A(n19471), .Y(n21174) );
  AOI222XL U23276 ( .A0(conv_3[287]), .A1(n16673), .B0(n22743), .B1(n21174), 
        .C0(conv_3[272]), .C1(n25289), .Y(n28276) );
  INVXL U23277 ( .A(n28276), .Y(n35139) );
  AOI22XL U23278 ( .A0(n16662), .A1(conv_3[392]), .B0(n25299), .B1(conv_3[362]), .Y(n18614) );
  NAND2XL U23279 ( .A(n18615), .B(n18614), .Y(n25716) );
  AOI22XL U23280 ( .A0(n25337), .A1(n35139), .B0(n25399), .B1(n25716), .Y(
        n18619) );
  INVXL U23281 ( .A(n25393), .Y(n25336) );
  INVXL U23282 ( .A(conv_3[422]), .Y(n30810) );
  AOI22XL U23283 ( .A0(n20735), .A1(conv_3[467]), .B0(conv_3[452]), .B1(n18634), .Y(n21172) );
  INVXL U23284 ( .A(conv_3[437]), .Y(n30816) );
  OAI222XL U23285 ( .A0(n30810), .A1(n22717), .B0(n22713), .B1(n21172), .C0(
        n19902), .C1(n30816), .Y(n28279) );
  AOI22XL U23286 ( .A0(n16662), .A1(conv_3[332]), .B0(n22690), .B1(conv_3[302]), .Y(n18616) );
  NAND2XL U23287 ( .A(n18617), .B(n18616), .Y(n25717) );
  AOI22XL U23288 ( .A0(n25336), .A1(n28279), .B0(n28289), .B1(n25717), .Y(
        n18618) );
  OAI211XL U23289 ( .A0(n35142), .A1(n16721), .B0(n18619), .C0(n18618), .Y(
        n26183) );
  AOI22XL U23290 ( .A0(n22762), .A1(conv_3[197]), .B0(n18240), .B1(conv_3[227]), .Y(n18621) );
  AOI22XL U23291 ( .A0(n16662), .A1(conv_3[212]), .B0(n22690), .B1(conv_3[182]), .Y(n18620) );
  NAND2XL U23292 ( .A(n18621), .B(n18620), .Y(n26182) );
  AOI22XL U23293 ( .A0(n25306), .A1(conv_3[137]), .B0(n22690), .B1(conv_3[122]), .Y(n18623) );
  NAND2XL U23294 ( .A(n18623), .B(n18622), .Y(n35140) );
  AOI22XL U23295 ( .A0(n22362), .A1(n26182), .B0(n28407), .B1(n35140), .Y(
        n18624) );
  NAND2XL U23296 ( .A(n16721), .B(n28278), .Y(n25720) );
  NAND2XL U23297 ( .A(n18624), .B(n25720), .Y(n25719) );
  AOI22XL U23298 ( .A0(n22762), .A1(conv_3[77]), .B0(n16673), .B1(conv_3[107]), 
        .Y(n18626) );
  AOI22XL U23299 ( .A0(n16662), .A1(conv_3[92]), .B0(n22690), .B1(conv_3[62]), 
        .Y(n18625) );
  NAND2XL U23300 ( .A(n18626), .B(n18625), .Y(n35148) );
  AOI22XL U23301 ( .A0(n22762), .A1(conv_3[17]), .B0(n25299), .B1(conv_3[2]), 
        .Y(n18628) );
  AOI22XL U23302 ( .A0(n16662), .A1(conv_3[32]), .B0(n18240), .B1(conv_3[47]), 
        .Y(n18627) );
  NAND2XL U23303 ( .A(n18628), .B(n18627), .Y(n28280) );
  AOI22XL U23304 ( .A0(n22362), .A1(n35148), .B0(n21100), .B1(n28280), .Y(
        n18629) );
  NAND2XL U23305 ( .A(n18629), .B(n25720), .Y(n25718) );
  AOI222XL U23306 ( .A0(n26183), .A1(n28467), .B0(n25719), .B1(n28465), .C0(
        n25718), .C1(n35130), .Y(n24567) );
  INVXL U23307 ( .A(n24567), .Y(n18650) );
  AOI22XL U23308 ( .A0(n16662), .A1(conv_3[331]), .B0(n18240), .B1(conv_3[346]), .Y(n18631) );
  AOI22XL U23309 ( .A0(n25306), .A1(conv_3[316]), .B0(n22690), .B1(conv_3[301]), .Y(n18630) );
  NAND2XL U23310 ( .A(n18631), .B(n18630), .Y(n25707) );
  INVXL U23311 ( .A(conv_3[466]), .Y(n30792) );
  AOI222XL U23312 ( .A0(n21144), .A1(n36246), .B0(n18658), .B1(conv_3[421]), 
        .C0(n21011), .C1(conv_3[436]), .Y(n25712) );
  AOI22XL U23313 ( .A0(n25306), .A1(conv_3[376]), .B0(n18240), .B1(conv_3[406]), .Y(n18633) );
  AOI22XL U23314 ( .A0(n16662), .A1(conv_3[391]), .B0(n22690), .B1(conv_3[361]), .Y(n18632) );
  NAND2XL U23315 ( .A(n18633), .B(n18632), .Y(n25715) );
  OAI2BB2XL U23316 ( .B0(n25712), .B1(n25393), .A0N(n25399), .A1N(n25715), .Y(
        n18636) );
  AOI22XL U23317 ( .A0(n20735), .A1(conv_3[526]), .B0(conv_3[511]), .B1(n18634), .Y(n21147) );
  AOI22XL U23318 ( .A0(n20735), .A1(conv_3[496]), .B0(conv_3[481]), .B1(n18634), .Y(n21148) );
  INVXL U23319 ( .A(n35153), .Y(n28301) );
  INVXL U23320 ( .A(conv_3[256]), .Y(n30597) );
  AOI222XL U23321 ( .A0(n21150), .A1(n21688), .B0(n16673), .B1(conv_3[286]), 
        .C0(conv_3[271]), .C1(n25289), .Y(n35157) );
  OAI22XL U23322 ( .A0(n28301), .A1(n16721), .B0(n35157), .B1(n25402), .Y(
        n18635) );
  AOI211XL U23323 ( .A0(n28289), .A1(n25707), .B0(n18636), .C0(n18635), .Y(
        n26177) );
  INVXL U23324 ( .A(n26177), .Y(n18648) );
  AOI22XL U23325 ( .A0(n16662), .A1(conv_3[211]), .B0(n18240), .B1(conv_3[226]), .Y(n18638) );
  AOI22XL U23326 ( .A0(n22762), .A1(conv_3[196]), .B0(n22690), .B1(conv_3[181]), .Y(n18637) );
  NAND2XL U23327 ( .A(n18638), .B(n18637), .Y(n35151) );
  AOI22XL U23328 ( .A0(n22762), .A1(conv_3[136]), .B0(n18810), .B1(conv_3[151]), .Y(n18640) );
  AOI22XL U23329 ( .A0(n18658), .A1(conv_3[121]), .B0(n18240), .B1(conv_3[166]), .Y(n18639) );
  NAND2XL U23330 ( .A(n18640), .B(n18639), .Y(n35154) );
  AOI22XL U23331 ( .A0(n22362), .A1(n35151), .B0(n21100), .B1(n35154), .Y(
        n18641) );
  NAND2XL U23332 ( .A(n16721), .B(n35153), .Y(n18646) );
  NAND2XL U23333 ( .A(n18641), .B(n18646), .Y(n25709) );
  AOI22XL U23334 ( .A0(n25306), .A1(conv_3[76]), .B0(n16662), .B1(conv_3[91]), 
        .Y(n18643) );
  AOI22XL U23335 ( .A0(n18658), .A1(conv_3[61]), .B0(n18240), .B1(conv_3[106]), 
        .Y(n18642) );
  NAND2XL U23336 ( .A(n18643), .B(n18642), .Y(n35152) );
  AOI22XL U23337 ( .A0(n25306), .A1(conv_3[16]), .B0(n22690), .B1(conv_3[1]), 
        .Y(n18645) );
  AOI22XL U23338 ( .A0(n16662), .A1(conv_3[31]), .B0(n18240), .B1(conv_3[46]), 
        .Y(n18644) );
  NAND2XL U23339 ( .A(n18645), .B(n18644), .Y(n26179) );
  AOI22XL U23340 ( .A0(n22362), .A1(n35152), .B0(n21100), .B1(n26179), .Y(
        n18647) );
  NAND2XL U23341 ( .A(n18647), .B(n18646), .Y(n25708) );
  AOI222XL U23342 ( .A0(n18648), .A1(n28467), .B0(n25709), .B1(n28465), .C0(
        n25708), .C1(n26470), .Y(n35017) );
  AOI222XL U23343 ( .A0(pool[115]), .A1(pool[116]), .B0(pool[115]), .B1(n35017), .C0(pool[116]), .C1(n35017), .Y(n18649) );
  AOI222XL U23344 ( .A0(n24568), .A1(n18650), .B0(n24568), .B1(n18649), .C0(
        n18650), .C1(n18649), .Y(n18651) );
  AOI222XL U23345 ( .A0(n35019), .A1(pool[118]), .B0(n35019), .B1(n18651), 
        .C0(pool[118]), .C1(n18651), .Y(n18652) );
  AOI22XL U23346 ( .A0(n16666), .A1(conv_3[209]), .B0(n16662), .B1(conv_3[224]), .Y(n18655) );
  NAND2XL U23347 ( .A(n18655), .B(n18654), .Y(n35167) );
  AOI22XL U23348 ( .A0(n20735), .A1(conv_3[539]), .B0(conv_3[524]), .B1(n19253), .Y(n21388) );
  AOI22XL U23349 ( .A0(n35269), .A1(conv_3[509]), .B0(conv_3[494]), .B1(n19253), .Y(n20538) );
  AOI22XL U23350 ( .A0(n16670), .A1(n35167), .B0(n35169), .B1(n28571), .Y(
        n18671) );
  INVX2 U23351 ( .A(n26621), .Y(n28366) );
  INVXL U23352 ( .A(conv_3[179]), .Y(n32226) );
  INVXL U23353 ( .A(conv_3[149]), .Y(n32175) );
  INVXL U23354 ( .A(conv_3[164]), .Y(n32256) );
  OAI22XL U23355 ( .A0(n19902), .A1(n32175), .B0(n22612), .B1(n32256), .Y(
        n18656) );
  AOI211XL U23356 ( .A0(conv_3[134]), .A1(n22759), .B0(n18657), .C0(n18656), 
        .Y(n35172) );
  INVXL U23357 ( .A(n35172), .Y(n28264) );
  AOI22XL U23358 ( .A0(n21011), .A1(conv_3[89]), .B0(n16662), .B1(conv_3[104]), 
        .Y(n18660) );
  AOI22XL U23359 ( .A0(n18658), .A1(conv_3[74]), .B0(n16673), .B1(conv_3[119]), 
        .Y(n18659) );
  NAND2XL U23360 ( .A(n18660), .B(n18659), .Y(n35168) );
  AOI22XL U23361 ( .A0(n28366), .A1(n28264), .B0(n18463), .B1(n35168), .Y(
        n18670) );
  AOI22XL U23362 ( .A0(n16666), .A1(conv_3[389]), .B0(n16716), .B1(conv_3[404]), .Y(n18662) );
  AOI22XL U23363 ( .A0(n18658), .A1(conv_3[374]), .B0(n16673), .B1(conv_3[419]), .Y(n18661) );
  NAND2XL U23364 ( .A(n18662), .B(n18661), .Y(n26166) );
  AOI22XL U23365 ( .A0(n16716), .A1(conv_3[44]), .B0(n22759), .B1(conv_3[14]), 
        .Y(n18664) );
  AOI22XL U23366 ( .A0(n16666), .A1(conv_3[29]), .B0(n16673), .B1(conv_3[59]), 
        .Y(n18663) );
  NAND2XL U23367 ( .A(n18664), .B(n18663), .Y(n28265) );
  INVXL U23368 ( .A(n28265), .Y(n35178) );
  INVXL U23369 ( .A(conv_3[479]), .Y(n32189) );
  INVXL U23370 ( .A(conv_3[464]), .Y(n32247) );
  AOI22XL U23371 ( .A0(n20735), .A1(n32189), .B0(n32247), .B1(n18526), .Y(
        n21381) );
  AOI222XL U23372 ( .A0(n21381), .A1(n36246), .B0(n22759), .B1(conv_3[434]), 
        .C0(n21011), .C1(conv_3[449]), .Y(n35171) );
  OAI22XL U23373 ( .A0(n35178), .A1(n35198), .B0(n35171), .B1(n34958), .Y(
        n18668) );
  INVXL U23374 ( .A(conv_3[269]), .Y(n33911) );
  INVXL U23375 ( .A(conv_3[254]), .Y(n29129) );
  AOI22XL U23376 ( .A0(n20735), .A1(n33911), .B0(n29129), .B1(n18516), .Y(
        n20541) );
  AOI222XL U23377 ( .A0(n20541), .A1(n22743), .B0(n16673), .B1(conv_3[299]), 
        .C0(conv_3[284]), .C1(n25289), .Y(n35170) );
  INVXL U23378 ( .A(conv_3[359]), .Y(n32135) );
  INVXL U23379 ( .A(conv_3[329]), .Y(n33287) );
  INVXL U23380 ( .A(conv_3[344]), .Y(n32219) );
  OAI22XL U23381 ( .A0(n19902), .A1(n33287), .B0(n22612), .B1(n32219), .Y(
        n18665) );
  AOI211XL U23382 ( .A0(conv_3[314]), .A1(n22616), .B0(n18666), .C0(n18665), 
        .Y(n26163) );
  OAI22XL U23383 ( .A0(n35170), .A1(n28575), .B0(n26163), .B1(n28479), .Y(
        n18667) );
  AOI211XL U23384 ( .A0(n16667), .A1(n26166), .B0(n18668), .C0(n18667), .Y(
        n18669) );
  NAND3XL U23385 ( .A(n18671), .B(n18670), .C(n18669), .Y(n18720) );
  INVXL U23386 ( .A(conv_3[403]), .Y(n34003) );
  INVXL U23387 ( .A(conv_3[373]), .Y(n32121) );
  OAI22XL U23388 ( .A0(n22612), .A1(n34003), .B0(n22717), .B1(n32121), .Y(
        n18673) );
  INVXL U23389 ( .A(conv_3[388]), .Y(n34142) );
  INVXL U23390 ( .A(conv_3[418]), .Y(n32190) );
  OAI22XL U23391 ( .A0(n22546), .A1(n34142), .B0(n18321), .B1(n32190), .Y(
        n18672) );
  INVXL U23392 ( .A(n26280), .Y(n24876) );
  AOI22XL U23393 ( .A0(n22616), .A1(conv_3[133]), .B0(n18240), .B1(conv_3[178]), .Y(n18675) );
  AOI22XL U23394 ( .A0(n16666), .A1(conv_3[148]), .B0(n16662), .B1(conv_3[163]), .Y(n18674) );
  NAND2XL U23395 ( .A(n18675), .B(n18674), .Y(n35189) );
  AOI22XL U23396 ( .A0(n16667), .A1(n24876), .B0(n28324), .B1(n35189), .Y(
        n18688) );
  INVX4 U23397 ( .A(n34981), .Y(n34963) );
  INVXL U23398 ( .A(conv_3[268]), .Y(n33905) );
  INVXL U23399 ( .A(conv_3[253]), .Y(n29123) );
  AOI22XL U23400 ( .A0(n20735), .A1(n33905), .B0(n29123), .B1(n18526), .Y(
        n21410) );
  AOI222XL U23401 ( .A0(n21410), .A1(n22743), .B0(n16673), .B1(conv_3[298]), 
        .C0(conv_3[283]), .C1(n16662), .Y(n35186) );
  INVXL U23402 ( .A(n35186), .Y(n28365) );
  AOI22XL U23403 ( .A0(n21011), .A1(conv_3[208]), .B0(n16673), .B1(conv_3[238]), .Y(n18677) );
  AOI22XL U23404 ( .A0(n16662), .A1(conv_3[223]), .B0(n22759), .B1(conv_3[193]), .Y(n18676) );
  NAND2XL U23405 ( .A(n18677), .B(n18676), .Y(n35185) );
  AOI22XL U23406 ( .A0(n16666), .A1(conv_3[328]), .B0(n22759), .B1(conv_3[313]), .Y(n18679) );
  NAND2XL U23407 ( .A(n18679), .B(n18678), .Y(n26275) );
  AOI22XL U23408 ( .A0(n35269), .A1(conv_3[538]), .B0(conv_3[523]), .B1(n18516), .Y(n20553) );
  AOI22XL U23409 ( .A0(n35269), .A1(conv_3[508]), .B0(conv_3[493]), .B1(n18526), .Y(n20554) );
  INVXL U23410 ( .A(n28364), .Y(n35183) );
  INVXL U23411 ( .A(conv_3[478]), .Y(n32326) );
  INVXL U23412 ( .A(conv_3[463]), .Y(n32241) );
  AOI22XL U23413 ( .A0(n35269), .A1(n32326), .B0(n32241), .B1(n18526), .Y(
        n21402) );
  AOI222XL U23414 ( .A0(n21402), .A1(n36246), .B0(n22690), .B1(conv_3[433]), 
        .C0(n22770), .C1(conv_3[448]), .Y(n35182) );
  OAI22XL U23415 ( .A0(n28551), .A1(n35183), .B0(n35182), .B1(n34958), .Y(
        n18685) );
  AOI22XL U23416 ( .A0(n16716), .A1(conv_3[43]), .B0(n22759), .B1(conv_3[13]), 
        .Y(n18681) );
  AOI22XL U23417 ( .A0(n22347), .A1(conv_3[28]), .B0(n16673), .B1(conv_3[58]), 
        .Y(n18680) );
  NAND2XL U23418 ( .A(n18681), .B(n18680), .Y(n35180) );
  INVXL U23419 ( .A(n35180), .Y(n28363) );
  AOI22XL U23420 ( .A0(n16662), .A1(conv_3[103]), .B0(n18658), .B1(conv_3[73]), 
        .Y(n18683) );
  AOI22XL U23421 ( .A0(n21011), .A1(conv_3[88]), .B0(n16673), .B1(conv_3[118]), 
        .Y(n18682) );
  NAND2XL U23422 ( .A(n18683), .B(n18682), .Y(n35179) );
  OAI2BB2XL U23423 ( .B0(n28363), .B1(n35198), .A0N(n35179), .A1N(n18463), .Y(
        n18684) );
  AOI211XL U23424 ( .A0(n34992), .A1(n26275), .B0(n18685), .C0(n18684), .Y(
        n18686) );
  NAND3XL U23425 ( .A(n18688), .B(n18687), .C(n18686), .Y(n18713) );
  AOI22XL U23426 ( .A0(n16662), .A1(conv_3[342]), .B0(n22759), .B1(conv_3[312]), .Y(n18690) );
  AOI22XL U23427 ( .A0(n16666), .A1(conv_3[327]), .B0(n18240), .B1(conv_3[357]), .Y(n18689) );
  NAND2XL U23428 ( .A(n18690), .B(n18689), .Y(n26259) );
  AOI22XL U23429 ( .A0(n21011), .A1(conv_3[27]), .B0(n16662), .B1(conv_3[42]), 
        .Y(n18692) );
  AOI22XL U23430 ( .A0(n22759), .A1(conv_3[12]), .B0(n16673), .B1(conv_3[57]), 
        .Y(n18691) );
  NAND2XL U23431 ( .A(n18692), .B(n18691), .Y(n28371) );
  AOI22XL U23432 ( .A0(n16659), .A1(n26259), .B0(n18197), .B1(n28371), .Y(
        n18705) );
  INVXL U23433 ( .A(conv_3[267]), .Y(n33479) );
  INVXL U23434 ( .A(conv_3[252]), .Y(n29182) );
  AOI22XL U23435 ( .A0(n35269), .A1(n33479), .B0(n29182), .B1(n19855), .Y(
        n21431) );
  AOI222XL U23436 ( .A0(n21431), .A1(n21688), .B0(n16673), .B1(conv_3[297]), 
        .C0(conv_3[282]), .C1(n16662), .Y(n35197) );
  INVXL U23437 ( .A(n35197), .Y(n28373) );
  AOI22XL U23438 ( .A0(n16662), .A1(conv_3[162]), .B0(n22690), .B1(conv_3[132]), .Y(n18694) );
  NAND2XL U23439 ( .A(n18694), .B(n18693), .Y(n35193) );
  AOI22XL U23440 ( .A0(n16662), .A1(conv_3[402]), .B0(n22690), .B1(conv_3[372]), .Y(n18696) );
  NAND2XL U23441 ( .A(n18696), .B(n18695), .Y(n26261) );
  INVXL U23442 ( .A(conv_3[477]), .Y(n32332) );
  INVXL U23443 ( .A(conv_3[462]), .Y(n31518) );
  AOI22XL U23444 ( .A0(n35269), .A1(n32332), .B0(n31518), .B1(n18516), .Y(
        n21423) );
  AOI222XL U23445 ( .A0(n21423), .A1(n36246), .B0(n18658), .B1(conv_3[432]), 
        .C0(n22770), .C1(conv_3[447]), .Y(n35201) );
  AOI2BB2XL U23446 ( .B0(n28556), .B1(n26261), .A0N(n34958), .A1N(n35201), .Y(
        n18703) );
  AOI22XL U23447 ( .A0(n35269), .A1(conv_3[537]), .B0(conv_3[522]), .B1(n19855), .Y(n19558) );
  AOI22XL U23448 ( .A0(n35269), .A1(conv_3[507]), .B0(conv_3[492]), .B1(n18634), .Y(n20563) );
  AOI22XL U23449 ( .A0(n22347), .A1(conv_3[207]), .B0(n16673), .B1(conv_3[237]), .Y(n18698) );
  AOI22XL U23450 ( .A0(n16662), .A1(conv_3[222]), .B0(n22690), .B1(conv_3[192]), .Y(n18697) );
  NAND2XL U23451 ( .A(n18698), .B(n18697), .Y(n28374) );
  INVXL U23452 ( .A(n28374), .Y(n35199) );
  AOI22XL U23453 ( .A0(n16662), .A1(conv_3[102]), .B0(n25299), .B1(conv_3[72]), 
        .Y(n18700) );
  AOI22XL U23454 ( .A0(n22347), .A1(conv_3[87]), .B0(n16673), .B1(conv_3[117]), 
        .Y(n18699) );
  NAND2XL U23455 ( .A(n18700), .B(n18699), .Y(n35194) );
  INVXL U23456 ( .A(n35194), .Y(n24881) );
  OAI22XL U23457 ( .A0(n35199), .A1(n28553), .B0(n24881), .B1(n16672), .Y(
        n18701) );
  AOI21XL U23458 ( .A0(n28571), .A1(n35206), .B0(n18701), .Y(n18702) );
  NAND4XL U23459 ( .A(n18705), .B(n18704), .C(n18703), .D(n18702), .Y(n18709)
         );
  NOR3XL U23460 ( .A(pool[119]), .B(n18713), .C(n18709), .Y(n18719) );
  NOR4BXL U23461 ( .AN(n18709), .B(n18708), .C(n18707), .D(n18706), .Y(n18715)
         );
  NAND2XL U23462 ( .A(pool[119]), .B(n18723), .Y(n18710) );
  NOR4BBXL U23463 ( .AN(n18713), .BN(n18712), .C(n18711), .D(n18710), .Y(
        n18714) );
  NAND4BBXL U23464 ( .AN(n18717), .BN(n18716), .C(n18715), .D(n18714), .Y(
        n18718) );
  OAI22XL U23465 ( .A0(n35018), .A1(pool[119]), .B0(n18723), .B1(n24569), .Y(
        n18724) );
  INVXL U23466 ( .A(n18724), .Y(N29335) );
  AOI22XL U23467 ( .A0(counter[3]), .A1(filter_1[53]), .B0(filter_1[5]), .B1(
        n20605), .Y(n18725) );
  AOI22XL U23468 ( .A0(n21011), .A1(pixel[49]), .B0(n18810), .B1(pixel[50]), 
        .Y(n18731) );
  AOI22XL U23469 ( .A0(n22759), .A1(pixel[48]), .B0(n16673), .B1(pixel[51]), 
        .Y(n18730) );
  AOI22XL U23470 ( .A0(n21011), .A1(pixel[45]), .B0(n18810), .B1(pixel[46]), 
        .Y(n18733) );
  AOI22XL U23471 ( .A0(n22759), .A1(pixel[44]), .B0(n16673), .B1(pixel[47]), 
        .Y(n18732) );
  AOI22XL U23472 ( .A0(n22369), .A1(n22171), .B0(n22370), .B1(n22169), .Y(
        n18739) );
  AOI22XL U23473 ( .A0(n21011), .A1(pixel[17]), .B0(n18810), .B1(pixel[18]), 
        .Y(n18735) );
  AOI22XL U23474 ( .A0(n22759), .A1(pixel[16]), .B0(n16673), .B1(pixel[19]), 
        .Y(n18734) );
  NAND2X1 U23475 ( .A(n18735), .B(n18734), .Y(n22170) );
  AOI22XL U23476 ( .A0(n18810), .A1(pixel[14]), .B0(n16673), .B1(pixel[15]), 
        .Y(n18737) );
  AOI22XL U23477 ( .A0(n21011), .A1(pixel[13]), .B0(n25299), .B1(pixel[12]), 
        .Y(n18736) );
  NAND2X1 U23478 ( .A(n18737), .B(n18736), .Y(n22172) );
  AOI22XL U23479 ( .A0(n22362), .A1(n22170), .B0(n21100), .B1(n22172), .Y(
        n18738) );
  AOI22XL U23480 ( .A0(n18810), .A1(pixel[26]), .B0(n25299), .B1(pixel[24]), 
        .Y(n18741) );
  AOI22XL U23481 ( .A0(n21011), .A1(pixel[25]), .B0(n16673), .B1(pixel[27]), 
        .Y(n18740) );
  AOI22XL U23482 ( .A0(n22616), .A1(pixel[56]), .B0(n16673), .B1(pixel[59]), 
        .Y(n18743) );
  AOI22XL U23483 ( .A0(n21011), .A1(pixel[57]), .B0(n18810), .B1(pixel[58]), 
        .Y(n18742) );
  AOI22XL U23484 ( .A0(pixel[55]), .A1(n16673), .B0(n25299), .B1(pixel[52]), 
        .Y(n18745) );
  AOI22XL U23485 ( .A0(n21011), .A1(pixel[53]), .B0(pixel[54]), .B1(n18810), 
        .Y(n18744) );
  AOI22XL U23486 ( .A0(n18810), .A1(pixel[22]), .B0(n25299), .B1(pixel[20]), 
        .Y(n18747) );
  AOI22XL U23487 ( .A0(n21011), .A1(pixel[21]), .B0(n16673), .B1(pixel[23]), 
        .Y(n18746) );
  NAND2X1 U23488 ( .A(n18747), .B(n18746), .Y(n22121) );
  AOI22XL U23489 ( .A0(n22370), .A1(n22122), .B0(n21100), .B1(n22121), .Y(
        n18748) );
  AOI22XL U23490 ( .A0(n16666), .A1(pixel[9]), .B0(n18810), .B1(pixel[10]), 
        .Y(n18752) );
  AOI22XL U23491 ( .A0(n22759), .A1(pixel[8]), .B0(n16673), .B1(pixel[11]), 
        .Y(n18751) );
  AOI22XL U23492 ( .A0(n18810), .A1(pixel[42]), .B0(n22616), .B1(pixel[40]), 
        .Y(n18754) );
  AOI22XL U23493 ( .A0(n20978), .A1(pixel[41]), .B0(n16673), .B1(pixel[43]), 
        .Y(n18753) );
  AOI22XL U23494 ( .A0(n21011), .A1(pixel[37]), .B0(n16673), .B1(pixel[39]), 
        .Y(n18756) );
  AOI22XL U23495 ( .A0(n18810), .A1(pixel[38]), .B0(n22616), .B1(pixel[36]), 
        .Y(n18755) );
  AOI22XL U23496 ( .A0(n21011), .A1(pixel[5]), .B0(n22616), .B1(pixel[4]), .Y(
        n18759) );
  AOI22XL U23497 ( .A0(n18810), .A1(pixel[6]), .B0(n16673), .B1(pixel[7]), .Y(
        n18758) );
  AOI22XL U23498 ( .A0(n26470), .A1(n23249), .B0(n16755), .B1(n22937), .Y(
        n18772) );
  AOI22XL U23499 ( .A0(n21011), .A1(pixel[1]), .B0(n16673), .B1(pixel[3]), .Y(
        n18763) );
  AOI22XL U23500 ( .A0(n22759), .A1(pixel[60]), .B0(n16673), .B1(pixel[63]), 
        .Y(n18765) );
  AOI22XL U23501 ( .A0(n21011), .A1(pixel[61]), .B0(n18810), .B1(pixel[62]), 
        .Y(n18764) );
  AOI22XL U23502 ( .A0(n21011), .A1(pixel[33]), .B0(n16673), .B1(pixel[35]), 
        .Y(n18767) );
  AOI22XL U23503 ( .A0(n18810), .A1(pixel[34]), .B0(n25299), .B1(pixel[32]), 
        .Y(n18766) );
  NAND2X1 U23504 ( .A(n18767), .B(n18766), .Y(n23239) );
  AOI22XL U23505 ( .A0(n21011), .A1(pixel[29]), .B0(n18810), .B1(pixel[30]), 
        .Y(n18769) );
  AOI22XL U23506 ( .A0(n22616), .A1(pixel[28]), .B0(n16673), .B1(pixel[31]), 
        .Y(n18768) );
  AOI22XL U23507 ( .A0(n22362), .A1(n23239), .B0(n21100), .B1(n23240), .Y(
        n18770) );
  OAI2BB1XL U23508 ( .A0N(n23252), .A1N(n18770), .B0(n16700), .Y(n18771) );
  AOI22XL U23509 ( .A0(n20978), .A1(pixel[6]), .B0(n18810), .B1(pixel[7]), .Y(
        n18775) );
  AOI22XL U23510 ( .A0(n22616), .A1(pixel[5]), .B0(n16673), .B1(pixel[8]), .Y(
        n18774) );
  NAND2X1 U23511 ( .A(n18775), .B(n18774), .Y(n22399) );
  AOI22XL U23512 ( .A0(n16666), .A1(pixel[2]), .B0(n22616), .B1(pixel[1]), .Y(
        n18779) );
  AOI22XL U23513 ( .A0(n16716), .A1(pixel[3]), .B0(n16723), .B1(pixel[4]), .Y(
        n18778) );
  NAND2X1 U23514 ( .A(n18779), .B(n18778), .Y(n22212) );
  AOI22XL U23515 ( .A0(n20978), .A1(pixel[34]), .B0(n18810), .B1(pixel[35]), 
        .Y(n18781) );
  AOI22XL U23516 ( .A0(n22616), .A1(pixel[33]), .B0(n16673), .B1(pixel[36]), 
        .Y(n18780) );
  NAND2X1 U23517 ( .A(n18781), .B(n18780), .Y(n22889) );
  AOI22XL U23518 ( .A0(n20978), .A1(pixel[38]), .B0(n18810), .B1(pixel[39]), 
        .Y(n18784) );
  AOI22XL U23519 ( .A0(n22616), .A1(pixel[37]), .B0(n16673), .B1(pixel[40]), 
        .Y(n18783) );
  NAND2X1 U23520 ( .A(n18784), .B(n18783), .Y(n22397) );
  AOI22XL U23521 ( .A0(n28366), .A1(n22889), .B0(n16670), .B1(n22397), .Y(
        n18785) );
  OAI2BB1XL U23522 ( .A0N(n26262), .A1N(n22212), .B0(n18785), .Y(n18819) );
  AOI22XL U23523 ( .A0(n16716), .A1(pixel[63]), .B0(n16673), .B1(pixel[0]), 
        .Y(n18787) );
  AOI22XL U23524 ( .A0(n21011), .A1(pixel[62]), .B0(n25299), .B1(pixel[61]), 
        .Y(n18786) );
  AOI22XL U23525 ( .A0(n20978), .A1(pixel[58]), .B0(n25299), .B1(pixel[57]), 
        .Y(n18789) );
  AOI22XL U23526 ( .A0(n18810), .A1(pixel[59]), .B0(n16673), .B1(pixel[60]), 
        .Y(n18788) );
  AOI22XL U23527 ( .A0(n20978), .A1(pixel[26]), .B0(n25299), .B1(pixel[25]), 
        .Y(n18791) );
  AOI22XL U23528 ( .A0(n18810), .A1(pixel[27]), .B0(n16673), .B1(pixel[28]), 
        .Y(n18790) );
  NAND2X1 U23529 ( .A(n18791), .B(n18790), .Y(n22202) );
  AOI22XL U23530 ( .A0(n22616), .A1(pixel[29]), .B0(n16673), .B1(pixel[32]), 
        .Y(n18793) );
  AOI22XL U23531 ( .A0(n21011), .A1(pixel[30]), .B0(n18810), .B1(pixel[31]), 
        .Y(n18792) );
  NAND2X1 U23532 ( .A(n18793), .B(n18792), .Y(n22210) );
  AOI22XL U23533 ( .A0(n18197), .A1(n22202), .B0(n18463), .B1(n22210), .Y(
        n18817) );
  AOI22XL U23534 ( .A0(n22616), .A1(pixel[21]), .B0(n16673), .B1(pixel[24]), 
        .Y(n18795) );
  AOI22XL U23535 ( .A0(n20978), .A1(pixel[22]), .B0(n18810), .B1(pixel[23]), 
        .Y(n18794) );
  NAND2X1 U23536 ( .A(n18795), .B(n18794), .Y(n22201) );
  AOI22XL U23537 ( .A0(n22616), .A1(pixel[49]), .B0(n16673), .B1(pixel[52]), 
        .Y(n18797) );
  AOI22XL U23538 ( .A0(n20978), .A1(pixel[50]), .B0(n18810), .B1(pixel[51]), 
        .Y(n18796) );
  AOI22XL U23539 ( .A0(n22362), .A1(n22201), .B0(n22370), .B1(n22396), .Y(
        n18803) );
  AOI22XL U23540 ( .A0(n20978), .A1(pixel[18]), .B0(n22616), .B1(pixel[17]), 
        .Y(n18799) );
  AOI22XL U23541 ( .A0(n16716), .A1(pixel[19]), .B0(n16723), .B1(pixel[20]), 
        .Y(n18798) );
  AOI22XL U23542 ( .A0(n22616), .A1(pixel[53]), .B0(n16673), .B1(pixel[56]), 
        .Y(n18801) );
  AOI22XL U23543 ( .A0(n20978), .A1(pixel[54]), .B0(n18810), .B1(pixel[55]), 
        .Y(n18800) );
  NAND2XL U23544 ( .A(n18801), .B(n18800), .Y(n22203) );
  AOI22XL U23545 ( .A0(n21100), .A1(n22402), .B0(n22369), .B1(n22203), .Y(
        n18802) );
  AOI22XL U23546 ( .A0(n20978), .A1(pixel[46]), .B0(n18810), .B1(pixel[47]), 
        .Y(n18805) );
  AOI22XL U23547 ( .A0(n22616), .A1(pixel[45]), .B0(n16723), .B1(pixel[48]), 
        .Y(n18804) );
  AOI22XL U23548 ( .A0(n22616), .A1(pixel[13]), .B0(n16673), .B1(pixel[16]), 
        .Y(n18807) );
  AOI22XL U23549 ( .A0(n20978), .A1(pixel[14]), .B0(n18810), .B1(pixel[15]), 
        .Y(n18806) );
  NAND2X1 U23550 ( .A(n18807), .B(n18806), .Y(n22845) );
  AOI22XL U23551 ( .A0(n18810), .A1(pixel[11]), .B0(n16673), .B1(pixel[12]), 
        .Y(n18809) );
  AOI22XL U23552 ( .A0(n20978), .A1(pixel[10]), .B0(n22616), .B1(pixel[9]), 
        .Y(n18808) );
  NAND2X1 U23553 ( .A(n18809), .B(n18808), .Y(n22843) );
  AOI22XL U23554 ( .A0(n22362), .A1(n22845), .B0(n21100), .B1(n22843), .Y(
        n18814) );
  AOI22XL U23555 ( .A0(n20978), .A1(pixel[42]), .B0(n18810), .B1(pixel[43]), 
        .Y(n18812) );
  AOI22XL U23556 ( .A0(n22616), .A1(pixel[41]), .B0(n16673), .B1(pixel[44]), 
        .Y(n18811) );
  NAND2XL U23557 ( .A(n22370), .B(n22846), .Y(n18813) );
  OAI211X1 U23558 ( .A0(n22401), .A1(n18815), .B0(n18814), .C0(n18813), .Y(
        n22818) );
  AOI22XL U23559 ( .A0(n34827), .A1(n22817), .B0(n16755), .B1(n22818), .Y(
        n18816) );
  OAI211XL U23560 ( .A0(n19143), .A1(n34989), .B0(n18817), .C0(n18816), .Y(
        n18818) );
  AOI211X4 U23561 ( .A0(n26376), .A1(n22399), .B0(n18819), .C0(n18818), .Y(
        n27860) );
  AOI22XL U23562 ( .A0(counter[3]), .A1(filter_1[52]), .B0(n20605), .B1(
        filter_1[4]), .Y(n18820) );
  OAI2BB1XL U23563 ( .A0N(n19004), .A1N(filter_1[34]), .B0(n18820), .Y(n18824)
         );
  AOI22XL U23564 ( .A0(n19006), .A1(filter_1[10]), .B0(n19005), .B1(
        filter_1[16]), .Y(n18823) );
  AOI22XL U23565 ( .A0(n19008), .A1(filter_1[46]), .B0(n19007), .B1(
        filter_1[28]), .Y(n18822) );
  AOI22XL U23566 ( .A0(n19009), .A1(filter_1[22]), .B0(n16676), .B1(
        filter_1[40]), .Y(n18821) );
  AOI22XL U23567 ( .A0(counter[3]), .A1(filter_1[51]), .B0(n19006), .B1(
        filter_1[9]), .Y(n18825) );
  OAI2BB1XL U23568 ( .A0N(n20605), .A1N(filter_1[3]), .B0(n18825), .Y(n18829)
         );
  AOI22XL U23569 ( .A0(n19008), .A1(filter_1[45]), .B0(n19005), .B1(
        filter_1[15]), .Y(n18828) );
  AOI22XL U23570 ( .A0(n19004), .A1(filter_1[33]), .B0(n16676), .B1(
        filter_1[39]), .Y(n18826) );
  INVXL U23571 ( .A(filter_1[20]), .Y(n28236) );
  AOI22XL U23572 ( .A0(n19008), .A1(filter_1[44]), .B0(n19005), .B1(
        filter_1[14]), .Y(n18830) );
  AOI22XL U23573 ( .A0(counter[3]), .A1(filter_1[48]), .B0(n20605), .B1(
        filter_1[0]), .Y(n18835) );
  NAND2XL U23574 ( .A(conv_1[465]), .B(n30672), .Y(n18847) );
  AOI22XL U23575 ( .A0(counter[3]), .A1(filter_1[49]), .B0(n16676), .B1(
        filter_1[37]), .Y(n18840) );
  OAI2BB1XL U23576 ( .A0N(n20605), .A1N(filter_1[1]), .B0(n18840), .Y(n18844)
         );
  AOI22XL U23577 ( .A0(n19004), .A1(filter_1[31]), .B0(n19007), .B1(
        filter_1[25]), .Y(n18843) );
  AOI22XL U23578 ( .A0(n19009), .A1(filter_1[19]), .B0(n19008), .B1(
        filter_1[43]), .Y(n18842) );
  AOI22XL U23579 ( .A0(n19006), .A1(filter_1[7]), .B0(n19005), .B1(
        filter_1[13]), .Y(n18841) );
  NAND2XL U23580 ( .A(n33507), .B(n27429), .Y(n18848) );
  INVXL U23581 ( .A(n18848), .Y(n18846) );
  AOI211XL U23582 ( .A0(n35272), .A1(n18847), .B0(n27860), .C0(n18846), .Y(
        n27013) );
  NAND2XL U23583 ( .A(n27013), .B(conv_1[466]), .Y(n27012) );
  NAND2XL U23584 ( .A(n18848), .B(n27012), .Y(n18850) );
  NAND2XL U23585 ( .A(n24909), .B(n18850), .Y(n18851) );
  NAND2XL U23586 ( .A(n33403), .B(n18850), .Y(n18849) );
  OAI31XL U23587 ( .A0(n33403), .A1(n27860), .A2(n18850), .B0(n18849), .Y(
        n26987) );
  NAND2XL U23588 ( .A(n26987), .B(conv_1[467]), .Y(n26986) );
  NOR2X1 U23589 ( .A(conv_1[472]), .B(n27602), .Y(n27601) );
  OAI21XL U23590 ( .A0(conv_1[473]), .A1(n27172), .B0(n32887), .Y(n26341) );
  INVXL U23591 ( .A(conv_1[474]), .Y(n26346) );
  INVXL U23592 ( .A(conv_1[470]), .Y(n20008) );
  NAND2XL U23593 ( .A(n27179), .B(conv_1[471]), .Y(n27603) );
  INVXL U23594 ( .A(conv_1[472]), .Y(n27604) );
  AOI21XL U23595 ( .A0(n32887), .A1(n29824), .B0(conv_1[476]), .Y(n29821) );
  INVXL U23596 ( .A(n29821), .Y(n29822) );
  NAND2XL U23597 ( .A(n32887), .B(n29824), .Y(n18858) );
  INVXL U23598 ( .A(conv_1[479]), .Y(n28738) );
  AND2X4 U23599 ( .A(ns[2]), .B(n20618), .Y(n29676) );
  INVXL U23600 ( .A(n18861), .Y(n18857) );
  AOI32XL U23601 ( .A0(n18858), .A1(n33506), .A2(n18857), .B0(n16658), .B1(
        n33506), .Y(n18859) );
  AOI21XL U23602 ( .A0(conv_1[476]), .A1(n18859), .B0(n35549), .Y(n18860) );
  OAI31XL U23603 ( .A0(n18861), .A1(n36001), .A2(n29822), .B0(n18860), .Y(
        n15987) );
  AOI22XL U23604 ( .A0(pixel[31]), .A1(n19475), .B0(pixel[29]), .B1(n16706), 
        .Y(n18865) );
  AOI22XL U23605 ( .A0(pixel[32]), .A1(n19099), .B0(pixel[27]), .B1(n21954), 
        .Y(n18864) );
  AOI22XL U23606 ( .A0(pixel[30]), .A1(n21887), .B0(pixel[28]), .B1(n16734), 
        .Y(n18863) );
  AOI22XL U23607 ( .A0(pixel[33]), .A1(n19097), .B0(pixel[34]), .B1(n19098), 
        .Y(n18862) );
  AOI22XL U23608 ( .A0(pixel[54]), .A1(n21887), .B0(pixel[58]), .B1(n19098), 
        .Y(n18868) );
  AOI22XL U23609 ( .A0(pixel[56]), .A1(n19099), .B0(pixel[52]), .B1(n16734), 
        .Y(n18867) );
  AOI22XL U23610 ( .A0(pixel[55]), .A1(n19475), .B0(pixel[57]), .B1(n19097), 
        .Y(n18866) );
  AOI22XL U23611 ( .A0(pixel[9]), .A1(n19097), .B0(pixel[10]), .B1(n19098), 
        .Y(n18873) );
  AOI22XL U23612 ( .A0(pixel[8]), .A1(n19099), .B0(pixel[4]), .B1(n16734), .Y(
        n18872) );
  AOI22XL U23613 ( .A0(pixel[5]), .A1(n22021), .B0(pixel[6]), .B1(n21887), .Y(
        n18871) );
  AOI22XL U23614 ( .A0(pixel[7]), .A1(n19475), .B0(pixel[3]), .B1(n21954), .Y(
        n18870) );
  AOI22XL U23615 ( .A0(pixel[62]), .A1(n21887), .B0(pixel[61]), .B1(n16706), 
        .Y(n18877) );
  AOI22XL U23616 ( .A0(pixel[60]), .A1(n16734), .B0(pixel[2]), .B1(n19098), 
        .Y(n18876) );
  AOI22XL U23617 ( .A0(pixel[0]), .A1(n19099), .B0(pixel[59]), .B1(n21954), 
        .Y(n18875) );
  AOI22XL U23618 ( .A0(pixel[63]), .A1(n19475), .B0(pixel[1]), .B1(n19097), 
        .Y(n18874) );
  INVXL U23619 ( .A(n23052), .Y(n23017) );
  AOI22XL U23620 ( .A0(pixel[38]), .A1(n21887), .B0(pixel[41]), .B1(n19097), 
        .Y(n18881) );
  AOI22XL U23621 ( .A0(pixel[40]), .A1(n19099), .B0(pixel[35]), .B1(n21954), 
        .Y(n18879) );
  AOI22XL U23622 ( .A0(pixel[39]), .A1(n19475), .B0(pixel[36]), .B1(n16734), 
        .Y(n18878) );
  AOI22XL U23623 ( .A0(pixel[49]), .A1(n19097), .B0(pixel[43]), .B1(n21954), 
        .Y(n18885) );
  AOI22XL U23624 ( .A0(pixel[50]), .A1(n19098), .B0(pixel[45]), .B1(n16706), 
        .Y(n18884) );
  AOI22XL U23625 ( .A0(pixel[44]), .A1(n16734), .B0(pixel[47]), .B1(n19475), 
        .Y(n18883) );
  AOI22XL U23626 ( .A0(pixel[48]), .A1(n19099), .B0(pixel[46]), .B1(n21887), 
        .Y(n18882) );
  AOI22XL U23627 ( .A0(pixel[21]), .A1(n22021), .B0(pixel[19]), .B1(n21954), 
        .Y(n18888) );
  AOI22XL U23628 ( .A0(pixel[15]), .A1(n19475), .B0(pixel[16]), .B1(n19099), 
        .Y(n18893) );
  AOI22XL U23629 ( .A0(pixel[14]), .A1(n21887), .B0(pixel[12]), .B1(n16734), 
        .Y(n18892) );
  AOI22XL U23630 ( .A0(pixel[17]), .A1(n19097), .B0(pixel[13]), .B1(n16706), 
        .Y(n18891) );
  AOI22XL U23631 ( .A0(pixel[18]), .A1(n19098), .B0(pixel[11]), .B1(n21954), 
        .Y(n18890) );
  AOI222XL U23632 ( .A0(n22450), .A1(n23278), .B0(n22153), .B1(n23276), .C0(
        n22449), .C1(n23272), .Y(n22265) );
  AOI22XL U23633 ( .A0(counter[3]), .A1(filter_2[53]), .B0(n19004), .B1(
        filter_2[35]), .Y(n18897) );
  AOI22XL U23634 ( .A0(counter[3]), .A1(filter_2[52]), .B0(n20605), .B1(
        filter_2[4]), .Y(n18902) );
  OAI2BB1XL U23635 ( .A0N(n16676), .A1N(filter_2[40]), .B0(n18902), .Y(n18906)
         );
  AOI22XL U23636 ( .A0(n19006), .A1(filter_2[10]), .B0(n19008), .B1(
        filter_2[46]), .Y(n18904) );
  AOI22XL U23637 ( .A0(n19009), .A1(filter_2[22]), .B0(n19004), .B1(
        filter_2[34]), .Y(n18903) );
  NAND2XL U23638 ( .A(n33424), .B(n29046), .Y(n18934) );
  INVXL U23639 ( .A(conv_2[498]), .Y(n34104) );
  AOI22XL U23640 ( .A0(counter[3]), .A1(filter_2[49]), .B0(n20605), .B1(
        filter_2[1]), .Y(n18907) );
  OAI2BB1XL U23641 ( .A0N(n19006), .A1N(filter_2[7]), .B0(n18907), .Y(n18911)
         );
  AOI22XL U23642 ( .A0(n19008), .A1(filter_2[43]), .B0(n19004), .B1(
        filter_2[31]), .Y(n18908) );
  INVX2 U23643 ( .A(n28126), .Y(n18913) );
  AOI22XL U23644 ( .A0(n19007), .A1(filter_2[24]), .B0(n20605), .B1(
        filter_2[0]), .Y(n18914) );
  INVX2 U23645 ( .A(n28124), .Y(n33989) );
  NAND2XL U23646 ( .A(n22883), .B(conv_2[495]), .Y(n22882) );
  OAI21XL U23647 ( .A0(n33422), .A1(n18913), .B0(n22882), .Y(n34232) );
  AOI22XL U23648 ( .A0(counter[3]), .A1(filter_2[50]), .B0(n20605), .B1(
        filter_2[2]), .Y(n18919) );
  OAI2BB1XL U23649 ( .A0N(n19009), .A1N(filter_2[20]), .B0(n18919), .Y(n18923)
         );
  NAND2XL U23650 ( .A(n33424), .B(n28128), .Y(n18924) );
  AOI22XL U23651 ( .A0(counter[3]), .A1(filter_2[51]), .B0(n20605), .B1(
        filter_2[3]), .Y(n18926) );
  OAI2BB1XL U23652 ( .A0N(n19008), .A1N(filter_2[45]), .B0(n18926), .Y(n18930)
         );
  AOI22XL U23653 ( .A0(n19009), .A1(filter_2[21]), .B0(n19006), .B1(
        filter_2[9]), .Y(n18927) );
  NAND2XL U23654 ( .A(n33424), .B(n28068), .Y(n18931) );
  NAND2XL U23655 ( .A(n18932), .B(n18931), .Y(n34100) );
  INVXL U23656 ( .A(n18941), .Y(n18937) );
  AOI32XL U23657 ( .A0(n18938), .A1(n36091), .A2(n18937), .B0(n16655), .B1(
        n36091), .Y(n18939) );
  AOI21XL U23658 ( .A0(conv_2[501]), .A1(n18939), .B0(n16651), .Y(n18940) );
  OAI31XL U23659 ( .A0(n18941), .A1(n34389), .A2(n30909), .B0(n18940), .Y(
        n14872) );
  INVXL U23660 ( .A(conv_2[275]), .Y(n28011) );
  NAND2X1 U23661 ( .A(n18945), .B(n18944), .Y(n22804) );
  AOI22XL U23662 ( .A0(n22362), .A1(n19051), .B0(n21100), .B1(n19050), .Y(
        n18947) );
  AOI22XL U23663 ( .A0(n22369), .A1(n23240), .B0(n22370), .B1(n22802), .Y(
        n18946) );
  AOI22XL U23664 ( .A0(n26470), .A1(n22804), .B0(n16755), .B1(n22123), .Y(
        n18951) );
  NAND2X1 U23665 ( .A(n18949), .B(n18948), .Y(n22803) );
  NAND2XL U23666 ( .A(n34827), .B(n22803), .Y(n18950) );
  INVX2 U23667 ( .A(n34711), .Y(n33994) );
  INVXL U23668 ( .A(conv_2[270]), .Y(n24041) );
  NOR4XL U23669 ( .A(n18913), .B(n33989), .C(n33994), .D(n24041), .Y(n18953)
         );
  NAND2XL U23670 ( .A(conv_2[270]), .B(n28124), .Y(n33993) );
  NAND2XL U23671 ( .A(n18913), .B(n33993), .Y(n18952) );
  OAI211XL U23672 ( .A0(n18913), .A1(n33993), .B0(n34711), .C0(n18952), .Y(
        n24552) );
  OR2XL U23673 ( .A(n18953), .B(n24550), .Y(n18954) );
  AOI21XL U23674 ( .A0(n28128), .A1(n34711), .B0(n18954), .Y(n23873) );
  INVXL U23675 ( .A(conv_2[272]), .Y(n23878) );
  NAND2XL U23676 ( .A(n28128), .B(n18954), .Y(n23874) );
  OAI21XL U23677 ( .A0(n23873), .A1(n23878), .B0(n23874), .Y(n23702) );
  AND2XL U23678 ( .A(n28883), .B(n18955), .Y(n28006) );
  INVXL U23679 ( .A(n28883), .Y(n35950) );
  INVXL U23680 ( .A(n28024), .Y(n28025) );
  AOI2BB1XL U23681 ( .A0N(n18956), .A1N(n28023), .B0(n16654), .Y(n18957) );
  INVXL U23682 ( .A(conv_2[284]), .Y(n28890) );
  AOI221XL U23683 ( .A0(n18957), .A1(conv_2[276]), .B0(n35952), .B1(
        conv_2[276]), .C0(n16651), .Y(n18958) );
  OAI31XL U23684 ( .A0(n28023), .A1(n16654), .A2(n28025), .B0(n18958), .Y(
        n15022) );
  AOI22XL U23685 ( .A0(n22370), .A1(n22121), .B0(n21100), .B1(n22122), .Y(
        n18959) );
  AND2X1 U23686 ( .A(n22936), .B(n16700), .Y(n18968) );
  AOI22XL U23687 ( .A0(n26263), .A1(n22170), .B0(n35195), .B1(n22169), .Y(
        n18966) );
  AOI22XL U23688 ( .A0(n28556), .A1(n22172), .B0(n35236), .B1(n22171), .Y(
        n18965) );
  INVX2 U23689 ( .A(n28277), .Y(n22847) );
  AOI22XL U23690 ( .A0(n34992), .A1(n23241), .B0(n35181), .B1(n23243), .Y(
        n18963) );
  NAND4X1 U23691 ( .A(n18966), .B(n18965), .C(n18964), .D(n18963), .Y(n18967)
         );
  INVXL U23692 ( .A(conv_2[66]), .Y(n30105) );
  INVXL U23693 ( .A(conv_2[64]), .Y(n25280) );
  NAND2XL U23694 ( .A(n29046), .B(n34699), .Y(n18970) );
  NAND2XL U23695 ( .A(conv_2[60]), .B(n23832), .Y(n23831) );
  OAI2BB1XL U23696 ( .A0N(n28126), .A1N(n34699), .B0(n23831), .Y(n35849) );
  AOI222XL U23697 ( .A0(n26742), .A1(n26743), .B0(n26742), .B1(conv_2[63]), 
        .C0(n26743), .C1(conv_2[63]), .Y(n18969) );
  NAND2XL U23698 ( .A(n18970), .B(n18969), .Y(n25276) );
  NAND2XL U23699 ( .A(n30242), .B(n18971), .Y(n30113) );
  NAND2XL U23700 ( .A(conv_2[65]), .B(n30113), .Y(n30101) );
  AOI221XL U23701 ( .A0(n30107), .A1(n18972), .B0(n33735), .B1(n18972), .C0(
        n36001), .Y(n18973) );
  AOI221XL U23702 ( .A0(n18973), .A1(conv_2[67]), .B0(n33730), .B1(conv_2[67]), 
        .C0(n16651), .Y(n18974) );
  OAI31XL U23703 ( .A0(n18975), .A1(n16654), .A2(n30106), .B0(n18974), .Y(
        n15161) );
  AOI22XL U23704 ( .A0(counter[3]), .A1(filter_3[53]), .B0(n19005), .B1(
        filter_3[17]), .Y(n18976) );
  AOI22XL U23705 ( .A0(counter[3]), .A1(filter_3[52]), .B0(n19005), .B1(
        filter_3[16]), .Y(n18981) );
  OAI2BB1XL U23706 ( .A0N(n20605), .A1N(filter_3[4]), .B0(n18981), .Y(n18985)
         );
  AOI22XL U23707 ( .A0(n19004), .A1(filter_3[34]), .B0(n16676), .B1(
        filter_3[40]), .Y(n18984) );
  AOI22XL U23708 ( .A0(n19009), .A1(filter_3[22]), .B0(n19008), .B1(
        filter_3[46]), .Y(n18983) );
  AOI22XL U23709 ( .A0(counter[3]), .A1(filter_3[51]), .B0(n20605), .B1(
        filter_3[3]), .Y(n18986) );
  OAI2BB1XL U23710 ( .A0N(n19008), .A1N(filter_3[45]), .B0(n18986), .Y(n18990)
         );
  NAND2XL U23711 ( .A(n29677), .B(n33509), .Y(n19018) );
  NAND2XL U23712 ( .A(filter_3[14]), .B(n19005), .Y(n18991) );
  AOI22XL U23713 ( .A0(counter[3]), .A1(filter_3[48]), .B0(n20605), .B1(
        filter_3[0]), .Y(n18998) );
  OAI2BB1XL U23714 ( .A0N(n19008), .A1N(filter_3[42]), .B0(n18998), .Y(n19002)
         );
  INVX2 U23715 ( .A(n29678), .Y(n27620) );
  NOR2X1 U23716 ( .A(n27620), .B(n27860), .Y(n31377) );
  NAND2XL U23717 ( .A(n31377), .B(conv_3[465]), .Y(n31376) );
  AOI22XL U23718 ( .A0(counter[3]), .A1(filter_3[49]), .B0(n20605), .B1(
        filter_3[1]), .Y(n19003) );
  OAI2BB1XL U23719 ( .A0N(n19004), .A1N(filter_3[31]), .B0(n19003), .Y(n19013)
         );
  AOI22XL U23720 ( .A0(n19006), .A1(filter_3[7]), .B0(n19005), .B1(
        filter_3[13]), .Y(n19012) );
  AOI22XL U23721 ( .A0(n19007), .A1(filter_3[25]), .B0(n16676), .B1(
        filter_3[37]), .Y(n19011) );
  AOI22XL U23722 ( .A0(n19009), .A1(filter_3[19]), .B0(n19008), .B1(
        filter_3[43]), .Y(n19010) );
  NAND2XL U23723 ( .A(n19015), .B(n29680), .Y(n19016) );
  NAND2XL U23724 ( .A(n30790), .B(conv_3[466]), .Y(n30789) );
  INVXL U23725 ( .A(conv_3[470]), .Y(n26124) );
  NAND2XL U23726 ( .A(n35810), .B(n32185), .Y(n19023) );
  NAND2BXL U23727 ( .AN(conv_3[475]), .B(n19023), .Y(n19026) );
  INVXL U23728 ( .A(n19027), .Y(n19022) );
  AOI32XL U23729 ( .A0(n19023), .A1(n35813), .A2(n19022), .B0(n16654), .B1(
        n35813), .Y(n19024) );
  AOI21XL U23730 ( .A0(conv_3[475]), .A1(n19024), .B0(n16653), .Y(n19025) );
  OAI31XL U23731 ( .A0(n19027), .A1(n36042), .A2(n19026), .B0(n19025), .Y(
        n15428) );
  AOI22XL U23732 ( .A0(n22362), .A1(n22204), .B0(n22369), .B1(n22202), .Y(
        n19031) );
  AOI22XL U23733 ( .A0(n22370), .A1(n22201), .B0(n21100), .B1(n22203), .Y(
        n19030) );
  AOI22XL U23734 ( .A0(n22370), .A1(n22397), .B0(n21100), .B1(n22399), .Y(
        n19033) );
  AOI22XL U23735 ( .A0(n22362), .A1(n22843), .B0(n22369), .B1(n22846), .Y(
        n19032) );
  NAND2X1 U23736 ( .A(n19033), .B(n19032), .Y(n23091) );
  AOI22XL U23737 ( .A0(n22362), .A1(n22402), .B0(n21100), .B1(n22845), .Y(
        n19035) );
  NAND2XL U23738 ( .A(n22369), .B(n22396), .Y(n19034) );
  AOI22XL U23739 ( .A0(n26470), .A1(n23091), .B0(n28465), .B1(n23092), .Y(
        n19036) );
  INVXL U23740 ( .A(n28161), .Y(n28191) );
  NAND4XL U23741 ( .A(conv_2[255]), .B(n28126), .C(n28124), .D(n34422), .Y(
        n19039) );
  NAND2XL U23742 ( .A(conv_2[255]), .B(n28124), .Y(n19038) );
  INVXL U23743 ( .A(n19038), .Y(n34420) );
  AOI221XL U23744 ( .A0(n18913), .A1(n19038), .B0(n28126), .B1(n34420), .C0(
        n28721), .Y(n29869) );
  NAND2XL U23745 ( .A(conv_2[256]), .B(n29869), .Y(n29868) );
  NAND2XL U23746 ( .A(n19039), .B(n29868), .Y(n19041) );
  NAND2XL U23747 ( .A(n35853), .B(n19041), .Y(n19040) );
  OAI31XL U23748 ( .A0(n35853), .A1(n28721), .A2(n19041), .B0(n19040), .Y(
        n27047) );
  NAND2XL U23749 ( .A(n19041), .B(n28128), .Y(n19042) );
  OAI2BB1XL U23750 ( .A0N(conv_2[257]), .A1N(n27047), .B0(n19042), .Y(n32983)
         );
  AND2XL U23751 ( .A(n28161), .B(n19043), .Y(n28178) );
  INVXL U23752 ( .A(n19049), .Y(n19045) );
  AOI32XL U23753 ( .A0(n19046), .A1(n34601), .A2(n19045), .B0(n16654), .B1(
        n34601), .Y(n19047) );
  AOI21XL U23754 ( .A0(conv_2[262]), .A1(n19047), .B0(n16651), .Y(n19048) );
  OAI31XL U23755 ( .A0(n19049), .A1(n16654), .A2(n28190), .B0(n19048), .Y(
        n15031) );
  AOI22XL U23756 ( .A0(n26376), .A1(n23244), .B0(n26262), .B1(n19052), .Y(
        n19057) );
  AOI22XL U23757 ( .A0(n18463), .A1(n23240), .B0(n28324), .B1(n23239), .Y(
        n19054) );
  AOI22XL U23758 ( .A0(n18197), .A1(n22802), .B0(n16670), .B1(n23242), .Y(
        n19053) );
  NAND2XL U23759 ( .A(conv_3[450]), .B(n29678), .Y(n19058) );
  NAND2XL U23760 ( .A(n28718), .B(n29680), .Y(n22443) );
  AOI21XL U23761 ( .A0(n30536), .A1(n19058), .B0(n27644), .Y(n22444) );
  NAND2XL U23762 ( .A(conv_3[451]), .B(n22444), .Y(n22441) );
  NAND2XL U23763 ( .A(n22443), .B(n22441), .Y(n19060) );
  NAND2XL U23764 ( .A(n18997), .B(n19060), .Y(n19059) );
  OAI31XL U23765 ( .A0(n18997), .A1(n27644), .A2(n19060), .B0(n19059), .Y(
        n30508) );
  NAND2XL U23766 ( .A(n19060), .B(n27619), .Y(n19061) );
  OAI2BB1XL U23767 ( .A0N(conv_3[452]), .A1N(n30508), .B0(n19061), .Y(n23048)
         );
  NAND2XL U23768 ( .A(n31517), .B(n19062), .Y(n35797) );
  NAND2XL U23769 ( .A(conv_3[455]), .B(n35797), .Y(n31508) );
  NAND2XL U23770 ( .A(n33780), .B(n31513), .Y(n19064) );
  NAND2BXL U23771 ( .AN(conv_3[460]), .B(n19064), .Y(n19067) );
  INVXL U23772 ( .A(n19068), .Y(n19063) );
  AOI32XL U23773 ( .A0(n19064), .A1(n35805), .A2(n19063), .B0(n16654), .B1(
        n35805), .Y(n19065) );
  AOI21XL U23774 ( .A0(conv_3[460]), .A1(n19065), .B0(n16653), .Y(n19066) );
  OAI31XL U23775 ( .A0(n19068), .A1(n34389), .A2(n19067), .B0(n19066), .Y(
        n15438) );
  AOI22XL U23776 ( .A0(pixel[54]), .A1(n19475), .B0(pixel[53]), .B1(n21887), 
        .Y(n19072) );
  AOI22XL U23777 ( .A0(pixel[55]), .A1(n19099), .B0(pixel[51]), .B1(n16734), 
        .Y(n19071) );
  AOI22XL U23778 ( .A0(pixel[56]), .A1(n19097), .B0(pixel[50]), .B1(n21954), 
        .Y(n19070) );
  INVXL U23779 ( .A(n23274), .Y(n19106) );
  AOI22XL U23780 ( .A0(pixel[49]), .A1(n19098), .B0(pixel[46]), .B1(n19475), 
        .Y(n19075) );
  AOI22XL U23781 ( .A0(pixel[48]), .A1(n19097), .B0(pixel[47]), .B1(n19099), 
        .Y(n19074) );
  AOI22XL U23782 ( .A0(pixel[21]), .A1(n21887), .B0(pixel[25]), .B1(n19098), 
        .Y(n19080) );
  AOI22XL U23783 ( .A0(pixel[19]), .A1(n16734), .B0(pixel[20]), .B1(n16706), 
        .Y(n19079) );
  AOI22XL U23784 ( .A0(pixel[22]), .A1(n19475), .B0(pixel[18]), .B1(n21954), 
        .Y(n19078) );
  AOI22XL U23785 ( .A0(pixel[23]), .A1(n19099), .B0(pixel[24]), .B1(n19097), 
        .Y(n19077) );
  NAND4XL U23786 ( .A(n19080), .B(n19079), .C(n19078), .D(n19077), .Y(n23277)
         );
  AOI22XL U23787 ( .A0(pixel[13]), .A1(n21887), .B0(pixel[11]), .B1(n16734), 
        .Y(n19084) );
  AOI22XL U23788 ( .A0(pixel[17]), .A1(n19098), .B0(pixel[10]), .B1(n21954), 
        .Y(n19083) );
  AOI22XL U23789 ( .A0(pixel[15]), .A1(n19099), .B0(pixel[12]), .B1(n16706), 
        .Y(n19082) );
  AOI22XL U23790 ( .A0(pixel[14]), .A1(n19475), .B0(pixel[16]), .B1(n19097), 
        .Y(n19081) );
  AOI22XL U23791 ( .A0(pixel[37]), .A1(n21887), .B0(pixel[40]), .B1(n19097), 
        .Y(n19088) );
  AOI22XL U23792 ( .A0(pixel[35]), .A1(n16734), .B0(pixel[41]), .B1(n19098), 
        .Y(n19087) );
  AOI22XL U23793 ( .A0(pixel[38]), .A1(n19475), .B0(pixel[36]), .B1(n16706), 
        .Y(n19086) );
  AOI22XL U23794 ( .A0(pixel[39]), .A1(n19099), .B0(pixel[34]), .B1(n21954), 
        .Y(n19085) );
  AOI22XL U23795 ( .A0(pixel[62]), .A1(n19475), .B0(pixel[59]), .B1(n16734), 
        .Y(n19092) );
  AOI22XL U23796 ( .A0(pixel[63]), .A1(n19099), .B0(pixel[60]), .B1(n16706), 
        .Y(n19091) );
  AOI22XL U23797 ( .A0(pixel[61]), .A1(n21887), .B0(pixel[1]), .B1(n19098), 
        .Y(n19090) );
  AOI22XL U23798 ( .A0(pixel[0]), .A1(n19097), .B0(pixel[58]), .B1(n21954), 
        .Y(n19089) );
  AOI22XL U23799 ( .A0(pixel[27]), .A1(n16734), .B0(pixel[28]), .B1(n16706), 
        .Y(n19096) );
  AOI22XL U23800 ( .A0(pixel[30]), .A1(n19475), .B0(pixel[33]), .B1(n19098), 
        .Y(n19095) );
  AOI22XL U23801 ( .A0(pixel[32]), .A1(n19097), .B0(pixel[29]), .B1(n21887), 
        .Y(n19094) );
  AOI22XL U23802 ( .A0(pixel[31]), .A1(n19099), .B0(pixel[26]), .B1(n21954), 
        .Y(n19093) );
  NAND4XL U23803 ( .A(n19096), .B(n19095), .C(n19094), .D(n19093), .Y(n23273)
         );
  AOI22XL U23804 ( .A0(n23272), .A1(n23275), .B0(n23278), .B1(n23273), .Y(
        n19105) );
  AOI22XL U23805 ( .A0(pixel[8]), .A1(n19097), .B0(pixel[4]), .B1(n16706), .Y(
        n19103) );
  AOI22XL U23806 ( .A0(pixel[9]), .A1(n19098), .B0(pixel[3]), .B1(n16734), .Y(
        n19102) );
  AOI22XL U23807 ( .A0(pixel[7]), .A1(n19099), .B0(pixel[2]), .B1(n21954), .Y(
        n19101) );
  AOI22XL U23808 ( .A0(pixel[5]), .A1(n21887), .B0(pixel[6]), .B1(n19475), .Y(
        n19100) );
  OR2XL U23809 ( .A(n24180), .B(n18913), .Y(n29782) );
  OAI21XL U23810 ( .A0(n18913), .A1(n19108), .B0(n24180), .Y(n29781) );
  NAND2XL U23811 ( .A(conv_2[301]), .B(n29781), .Y(n19109) );
  OAI21XL U23812 ( .A0(n35853), .A1(n19108), .B0(n19110), .Y(n33057) );
  INVXL U23813 ( .A(n19111), .Y(n19112) );
  INVXL U23814 ( .A(conv_2[305]), .Y(n30861) );
  NAND2XL U23815 ( .A(n28918), .B(conv_2[306]), .Y(n28899) );
  INVXL U23816 ( .A(conv_2[307]), .Y(n28903) );
  NAND2XL U23817 ( .A(n29947), .B(conv_2[308]), .Y(n35969) );
  INVXL U23818 ( .A(conv_2[314]), .Y(n33985) );
  INVXL U23819 ( .A(n19119), .Y(n19115) );
  AOI32XL U23820 ( .A0(n19116), .A1(n35976), .A2(n19115), .B0(n36042), .B1(
        n35976), .Y(n19117) );
  AOI21XL U23821 ( .A0(conv_2[310]), .A1(n19117), .B0(n16651), .Y(n19118) );
  OAI31XL U23822 ( .A0(n19119), .A1(n16654), .A2(n28628), .B0(n19118), .Y(
        n14998) );
  INVXL U23823 ( .A(n22450), .Y(n19124) );
  AOI22XL U23824 ( .A0(n23783), .A1(n22266), .B0(n23785), .B1(n22449), .Y(
        n19123) );
  AOI22XL U23825 ( .A0(n23278), .A1(n22151), .B0(n23276), .B1(n22447), .Y(
        n19120) );
  INVXL U23826 ( .A(conv_1[140]), .Y(n26776) );
  NAND2XL U23827 ( .A(n27230), .B(n34740), .Y(n19131) );
  NAND2XL U23828 ( .A(n27429), .B(n34740), .Y(n19125) );
  NAND2XL U23829 ( .A(conv_1[135]), .B(n30672), .Y(n33501) );
  NAND2XL U23830 ( .A(n35272), .B(n33501), .Y(n19126) );
  OAI211XL U23831 ( .A0(n35272), .A1(n33501), .B0(n34740), .C0(n19126), .Y(
        n23943) );
  INVXL U23832 ( .A(conv_1[136]), .Y(n23945) );
  OAI21XL U23833 ( .A0(n33403), .A1(n34426), .B0(n19128), .Y(n19129) );
  INVXL U23834 ( .A(n19129), .Y(n26916) );
  AOI222XL U23835 ( .A0(n26749), .A1(n26748), .B0(n26749), .B1(conv_1[138]), 
        .C0(n26748), .C1(conv_1[138]), .Y(n19130) );
  AND2XL U23836 ( .A(n19131), .B(n19130), .Y(n26928) );
  NAND2XL U23837 ( .A(n35339), .B(n19132), .Y(n26771) );
  NAND2XL U23838 ( .A(n26776), .B(n26771), .Y(n26760) );
  INVXL U23839 ( .A(n35339), .Y(n32780) );
  OR2XL U23840 ( .A(n35339), .B(n19132), .Y(n26772) );
  AOI21XL U23841 ( .A0(conv_1[140]), .A1(n26772), .B0(n35339), .Y(n26759) );
  INVXL U23842 ( .A(conv_1[141]), .Y(n26764) );
  AOI21XL U23843 ( .A0(n35338), .A1(conv_1[142]), .B0(n35339), .Y(n26766) );
  INVXL U23844 ( .A(conv_1[145]), .Y(n19918) );
  NAND2XL U23845 ( .A(n35339), .B(n26754), .Y(n19134) );
  NAND2XL U23846 ( .A(n19918), .B(n19134), .Y(n19137) );
  INVXL U23847 ( .A(conv_1[149]), .Y(n26831) );
  INVXL U23848 ( .A(n19138), .Y(n19133) );
  AOI32XL U23849 ( .A0(n19134), .A1(n34271), .A2(n19133), .B0(n16655), .B1(
        n34271), .Y(n19135) );
  AOI21XL U23850 ( .A0(conv_1[145]), .A1(n19135), .B0(n35549), .Y(n19136) );
  OAI31XL U23851 ( .A0(n19138), .A1(n16654), .A2(n19137), .B0(n19136), .Y(
        n16318) );
  NAND2XL U23852 ( .A(n22362), .B(n22399), .Y(n19139) );
  AOI22XL U23853 ( .A0(n28366), .A1(n22202), .B0(n16670), .B1(n22210), .Y(
        n19142) );
  AOI22XL U23854 ( .A0(n35130), .A1(n22817), .B0(n34827), .B1(n22818), .Y(
        n19141) );
  AOI21X1 U23855 ( .A0(n16755), .A1(n22850), .B0(n19144), .Y(n19145) );
  BUFX4 U23856 ( .A(n19145), .Y(n27532) );
  INVXL U23857 ( .A(conv_1[384]), .Y(n34340) );
  NOR2X1 U23858 ( .A(n33423), .B(n27532), .Y(n23817) );
  NAND2X1 U23859 ( .A(n23817), .B(conv_1[375]), .Y(n23816) );
  INVXL U23860 ( .A(n23816), .Y(n19146) );
  AOI32XL U23861 ( .A0(n27535), .A1(n23816), .A2(n27429), .B0(n35272), .B1(
        n19146), .Y(n23822) );
  INVXL U23862 ( .A(conv_1[376]), .Y(n23824) );
  NOR2X1 U23863 ( .A(n19149), .B(n19148), .Y(n23724) );
  INVXL U23864 ( .A(n19150), .Y(n19151) );
  NOR2X1 U23865 ( .A(conv_1[380]), .B(n33177), .Y(n33176) );
  OAI21XL U23866 ( .A0(conv_1[383]), .A1(n35461), .B0(n35463), .Y(n34335) );
  NAND2XL U23867 ( .A(n23135), .B(conv_1[381]), .Y(n23129) );
  INVXL U23868 ( .A(conv_1[382]), .Y(n23133) );
  AOI21XL U23869 ( .A0(n35463), .A1(n33089), .B0(conv_1[386]), .Y(n33086) );
  INVXL U23870 ( .A(n33086), .Y(n33087) );
  NAND2XL U23871 ( .A(n35463), .B(n33089), .Y(n19155) );
  INVXL U23872 ( .A(conv_1[389]), .Y(n33152) );
  INVXL U23873 ( .A(n19158), .Y(n19154) );
  AOI32XL U23874 ( .A0(n19155), .A1(n35466), .A2(n19154), .B0(n16655), .B1(
        n35466), .Y(n19156) );
  AOI21XL U23875 ( .A0(conv_1[386]), .A1(n19156), .B0(n35549), .Y(n19157) );
  OAI31XL U23876 ( .A0(n19158), .A1(n36042), .A2(n33087), .B0(n19157), .Y(
        n16077) );
  AOI22XL U23877 ( .A0(n28414), .A1(n23241), .B0(n35181), .B1(n22169), .Y(
        n19162) );
  AOI22XL U23878 ( .A0(n28556), .A1(n22170), .B0(n22847), .B1(n23243), .Y(
        n19160) );
  AOI22XL U23879 ( .A0(n26263), .A1(n22121), .B0(n35195), .B1(n22171), .Y(
        n19159) );
  AND4X2 U23880 ( .A(n19162), .B(n19161), .C(n19160), .D(n19159), .Y(n19164)
         );
  NAND2XL U23881 ( .A(conv_2[90]), .B(n28124), .Y(n19166) );
  NAND2XL U23882 ( .A(n34448), .B(n28126), .Y(n19167) );
  INVXL U23883 ( .A(n19167), .Y(n19165) );
  AOI211XL U23884 ( .A0(n18913), .A1(n19166), .B0(n26509), .C0(n19165), .Y(
        n24483) );
  NAND2XL U23885 ( .A(conv_2[91]), .B(n24483), .Y(n24482) );
  NAND2XL U23886 ( .A(n19167), .B(n24482), .Y(n19169) );
  NAND2XL U23887 ( .A(n35853), .B(n19169), .Y(n19168) );
  OAI31XL U23888 ( .A0(n35853), .A1(n26509), .A2(n19169), .B0(n19168), .Y(
        n30007) );
  NAND2XL U23889 ( .A(n19169), .B(n28128), .Y(n19170) );
  OAI2BB1XL U23890 ( .A0N(conv_2[92]), .A1N(n30007), .B0(n19170), .Y(n23031)
         );
  NAND2XL U23891 ( .A(n30225), .B(n19171), .Y(n28691) );
  NAND2XL U23892 ( .A(conv_2[95]), .B(n28691), .Y(n28696) );
  INVXL U23893 ( .A(conv_2[96]), .Y(n19173) );
  NAND2XL U23894 ( .A(n19172), .B(n28690), .Y(n28694) );
  NAND2XL U23895 ( .A(n30940), .B(n28694), .Y(n28698) );
  NAND2XL U23896 ( .A(n19173), .B(n28698), .Y(n28701) );
  NAND2XL U23897 ( .A(n30940), .B(n28701), .Y(n19175) );
  INVXL U23898 ( .A(n19178), .Y(n19174) );
  AOI32XL U23899 ( .A0(n19175), .A1(n34447), .A2(n19174), .B0(n16655), .B1(
        n34447), .Y(n19176) );
  AOI21XL U23900 ( .A0(conv_2[97]), .A1(n19176), .B0(n16651), .Y(n19177) );
  OAI31XL U23901 ( .A0(n19178), .A1(n16654), .A2(n30203), .B0(n19177), .Y(
        n15141) );
  INVXL U23902 ( .A(n19244), .Y(n36249) );
  INVXL U23903 ( .A(n19179), .Y(n26039) );
  NAND2XL U23904 ( .A(n36245), .B(n16668), .Y(n35262) );
  INVXL U23905 ( .A(n35265), .Y(n19224) );
  NOR4XL U23906 ( .A(N18471), .B(cursor[6]), .C(n22612), .D(n19181), .Y(n35259) );
  NAND2XL U23907 ( .A(n21764), .B(n19182), .Y(n35260) );
  INVXL U23908 ( .A(conv_3[380]), .Y(n31459) );
  NAND2XL U23909 ( .A(conv_3[375]), .B(n29678), .Y(n27531) );
  NAND2XL U23910 ( .A(n29680), .B(n27535), .Y(n19188) );
  AOI211XL U23911 ( .A0(n30536), .A1(n27531), .B0(n27532), .C0(n19189), .Y(
        n30637) );
  INVXL U23912 ( .A(n19189), .Y(n19190) );
  OAI2BB1XL U23913 ( .A0N(conv_3[376]), .A1N(n30637), .B0(n19190), .Y(n24246)
         );
  AND2XL U23914 ( .A(n19192), .B(n19191), .Y(n24202) );
  NAND2XL U23915 ( .A(n34164), .B(n19194), .Y(n19195) );
  NAND2BXL U23916 ( .AN(conv_3[382]), .B(n19195), .Y(n31385) );
  INVXL U23917 ( .A(n19198), .Y(n31386) );
  INVXL U23918 ( .A(conv_3[389]), .Y(n32204) );
  AOI32XL U23919 ( .A0(n31386), .A1(n34168), .A2(n19195), .B0(n16658), .B1(
        n34168), .Y(n19196) );
  AOI21XL U23920 ( .A0(conv_3[382]), .A1(n19196), .B0(n31384), .Y(n19197) );
  OAI31XL U23921 ( .A0(n19198), .A1(n16658), .A2(n31385), .B0(n19197), .Y(
        n15491) );
  AOI222X1 U23922 ( .A0(n22448), .A1(n23278), .B0(n22449), .B1(n23276), .C0(
        n22447), .C1(n23272), .Y(n22157) );
  AOI22XL U23923 ( .A0(n34906), .A1(n22450), .B0(n23017), .B1(n22151), .Y(
        n19200) );
  AOI22XL U23924 ( .A0(n25766), .A1(n22152), .B0(n34921), .B1(n22266), .Y(
        n19199) );
  NAND4XL U23925 ( .A(conv_3[405]), .B(n29680), .C(n29678), .D(n34229), .Y(
        n19203) );
  NAND2XL U23926 ( .A(conv_3[405]), .B(n29678), .Y(n19202) );
  INVXL U23927 ( .A(n19202), .Y(n34228) );
  AOI221XL U23928 ( .A0(n30536), .A1(n19202), .B0(n29680), .B1(n34228), .C0(
        n28070), .Y(n30633) );
  NAND2XL U23929 ( .A(conv_3[406]), .B(n30633), .Y(n30632) );
  AND2XL U23930 ( .A(n19203), .B(n30632), .Y(n19204) );
  NAND2XL U23931 ( .A(n27619), .B(n34229), .Y(n19205) );
  AND2XL U23932 ( .A(n19205), .B(n19204), .Y(n30544) );
  AOI222XL U23933 ( .A0(n26814), .A1(n26815), .B0(n26814), .B1(conv_3[409]), 
        .C0(n26815), .C1(conv_3[409]), .Y(n19206) );
  AND2XL U23934 ( .A(n32558), .B(n19206), .Y(n32626) );
  AOI21XL U23935 ( .A0(conv_3[411]), .A1(n32005), .B0(n32557), .Y(n31987) );
  INVXL U23936 ( .A(conv_3[412]), .Y(n31992) );
  OAI21XL U23937 ( .A0(conv_3[411]), .A1(n32004), .B0(n32557), .Y(n31988) );
  NAND2XL U23938 ( .A(n32555), .B(n32556), .Y(n31993) );
  INVXL U23939 ( .A(conv_3[419]), .Y(n32196) );
  INVXL U23940 ( .A(n19211), .Y(n19208) );
  AOI32XL U23941 ( .A0(n32556), .A1(n34227), .A2(n19208), .B0(n16655), .B1(
        n34227), .Y(n19209) );
  AOI21XL U23942 ( .A0(conv_3[414]), .A1(n19209), .B0(n16653), .Y(n19210) );
  OAI31XL U23943 ( .A0(n19211), .A1(n16658), .A2(n31993), .B0(n19210), .Y(
        n15469) );
  INVXL U23944 ( .A(conv_1[300]), .Y(n33866) );
  NAND2XL U23945 ( .A(n33867), .B(n19213), .Y(n33864) );
  INVXL U23946 ( .A(n19214), .Y(n19212) );
  OAI211XL U23947 ( .A0(n19213), .A1(n27429), .B0(n33867), .C0(n19212), .Y(
        n24527) );
  INVXL U23948 ( .A(conv_1[301]), .Y(n24529) );
  NOR2X1 U23949 ( .A(n24527), .B(n24529), .Y(n24525) );
  OAI21XL U23950 ( .A0(n33403), .A1(n19108), .B0(n19215), .Y(n24515) );
  AOI21XL U23951 ( .A0(conv_1[302]), .A1(n24515), .B0(n24514), .Y(n19216) );
  NAND2XL U23952 ( .A(n27231), .B(n33867), .Y(n19217) );
  AND2XL U23953 ( .A(n19217), .B(n19216), .Y(n24225) );
  AOI21XL U23954 ( .A0(n24153), .A1(conv_1[306]), .B0(n28644), .Y(n22319) );
  INVXL U23955 ( .A(n28644), .Y(n24159) );
  AOI2BB1XL U23956 ( .A0N(n22319), .A1N(n19218), .B0(n16658), .Y(n19219) );
  INVXL U23957 ( .A(conv_1[314]), .Y(n24814) );
  AOI221XL U23958 ( .A0(n19219), .A1(conv_1[307]), .B0(n24151), .B1(
        conv_1[307]), .C0(n35549), .Y(n19220) );
  OAI31XL U23959 ( .A0(n22319), .A1(n16658), .A2(n22317), .B0(n19220), .Y(
        n16156) );
  AND2XL U23960 ( .A(n19221), .B(n35262), .Y(n19225) );
  NAND2XL U23961 ( .A(counter[2]), .B(n19245), .Y(n20163) );
  AOI21XL U23962 ( .A0(n19227), .A1(n20163), .B0(n19242), .Y(N30141) );
  NOR3XL U23963 ( .A(n19229), .B(n19228), .C(n19242), .Y(N30140) );
  AOI22XL U23964 ( .A0(n35265), .A1(n35258), .B0(n35256), .B1(add_x_358_n1), 
        .Y(n19230) );
  NAND2XL U23965 ( .A(cursor[6]), .B(n19230), .Y(n19231) );
  OAI22XL U23966 ( .A0(n19231), .A1(n35268), .B0(cursor[6]), .B1(n19230), .Y(
        n16644) );
  INVXL U23967 ( .A(pixel[8]), .Y(n19232) );
  INVXL U23968 ( .A(pixel[7]), .Y(n19233) );
  AOI22XL U23969 ( .A0(n22896), .A1(n19232), .B0(n19233), .B1(n23672), .Y(
        N17501) );
  INVXL U23970 ( .A(pixel[9]), .Y(n19234) );
  AOI22XL U23971 ( .A0(n22896), .A1(n19234), .B0(n19232), .B1(n23672), .Y(
        N17502) );
  INVXL U23972 ( .A(pixel[6]), .Y(n19239) );
  AOI22XL U23973 ( .A0(n22896), .A1(n19233), .B0(n19239), .B1(n23672), .Y(
        N17500) );
  INVXL U23974 ( .A(pixel[3]), .Y(n19236) );
  INVXL U23975 ( .A(pixel[2]), .Y(n20721) );
  AOI22XL U23976 ( .A0(n22896), .A1(n19236), .B0(n20721), .B1(n23672), .Y(
        N17496) );
  INVXL U23977 ( .A(pixel[11]), .Y(n23673) );
  INVXL U23978 ( .A(pixel[10]), .Y(n19235) );
  AOI22XL U23979 ( .A0(n22896), .A1(n23673), .B0(n19235), .B1(n23672), .Y(
        N17504) );
  AOI22XL U23980 ( .A0(n22896), .A1(n19235), .B0(n19234), .B1(n23672), .Y(
        N17503) );
  INVXL U23981 ( .A(pixel[5]), .Y(n19238) );
  INVXL U23982 ( .A(pixel[4]), .Y(n19237) );
  AOI22XL U23983 ( .A0(n22896), .A1(n19238), .B0(n19237), .B1(n23672), .Y(
        N17498) );
  AOI22XL U23984 ( .A0(n22896), .A1(n19237), .B0(n19236), .B1(n23672), .Y(
        N17497) );
  AOI22XL U23985 ( .A0(n22896), .A1(n19239), .B0(n19238), .B1(n23672), .Y(
        N17499) );
  NAND2X1 U23986 ( .A(n19243), .B(n19244), .Y(n33367) );
  INVXL U23987 ( .A(n33367), .Y(n19241) );
  OAI22XL U23988 ( .A0(counter[0]), .A1(n19242), .B0(n19241), .B1(n19240), .Y(
        n16636) );
  NAND3XL U23989 ( .A(n19247), .B(n19246), .C(n19245), .Y(n20599) );
  INVXL U23990 ( .A(weight_1_bias_3[0]), .Y(n19248) );
  NAND2XL U23991 ( .A(in_data[8]), .B(in_data[7]), .Y(n20168) );
  OAI22XL U23992 ( .A0(n36155), .A1(n19248), .B0(n36124), .B1(n36153), .Y(
        n14105) );
  INVXL U23993 ( .A(weight_1_bias_2[0]), .Y(n36138) );
  OAI22XL U23994 ( .A0(n36155), .A1(n36138), .B0(n36153), .B1(n19248), .Y(
        n14104) );
  OR2X1 U23995 ( .A(n36246), .B(n25123), .Y(n22014) );
  INVXL U23996 ( .A(conv_3[465]), .Y(n31379) );
  AOI2BB2X1 U23997 ( .B0(n20735), .B1(n31379), .A0N(conv_3[450]), .A1N(n35269), 
        .Y(n34951) );
  AOI22XL U23998 ( .A0(n21990), .A1(conv_3[420]), .B0(n21991), .B1(n34951), 
        .Y(n19252) );
  AOI22XL U23999 ( .A0(n21887), .A1(conv_3[435]), .B0(n21954), .B1(conv_3[390]), .Y(n19251) );
  AOI22XL U24000 ( .A0(n16734), .A1(conv_3[405]), .B0(n22015), .B1(conv_3[15]), 
        .Y(n19250) );
  NAND2XL U24001 ( .A(n21992), .B(conv_3[0]), .Y(n19249) );
  NAND4XL U24002 ( .A(n19252), .B(n19251), .C(n19250), .D(n19249), .Y(n34972)
         );
  AOI22XL U24003 ( .A0(n20735), .A1(conv_3[495]), .B0(conv_3[480]), .B1(n19253), .Y(n22226) );
  AOI22XL U24004 ( .A0(n20735), .A1(conv_3[525]), .B0(conv_3[510]), .B1(n19253), .Y(n22227) );
  INVXL U24005 ( .A(n34953), .Y(n21113) );
  INVXL U24006 ( .A(n25987), .Y(n26066) );
  INVXL U24007 ( .A(n22226), .Y(n34949) );
  AOI22XL U24008 ( .A0(n26066), .A1(n34949), .B0(n34903), .B1(n34951), .Y(
        n19259) );
  AOI22XL U24009 ( .A0(n20978), .A1(conv_3[105]), .B0(n22690), .B1(conv_3[90]), 
        .Y(n19254) );
  NAND2XL U24010 ( .A(n19255), .B(n19254), .Y(n34965) );
  AOI22XL U24011 ( .A0(n16666), .A1(conv_3[345]), .B0(n22616), .B1(conv_3[330]), .Y(n19257) );
  NAND2XL U24012 ( .A(n19257), .B(n19256), .Y(n34964) );
  AOI22XL U24013 ( .A0(n35236), .A1(n34965), .B0(n19179), .B1(n34964), .Y(
        n19258) );
  OAI211XL U24014 ( .A0(n21113), .A1(n23053), .B0(n19259), .C0(n19258), .Y(
        n19269) );
  INVXL U24015 ( .A(conv_3[255]), .Y(n30609) );
  INVXL U24016 ( .A(conv_3[240]), .Y(n30605) );
  AOI22XL U24017 ( .A0(n20735), .A1(n30609), .B0(n30605), .B1(n19253), .Y(
        n22235) );
  AOI22XL U24018 ( .A0(n21831), .A1(n22235), .B0(n34953), .B1(n21830), .Y(
        n34968) );
  AOI22XL U24019 ( .A0(n16666), .A1(conv_3[45]), .B0(n18240), .B1(conv_3[75]), 
        .Y(n19260) );
  NAND2XL U24020 ( .A(n19261), .B(n19260), .Y(n34962) );
  AOI222XL U24021 ( .A0(n22235), .A1(n36246), .B0(n18658), .B1(conv_3[210]), 
        .C0(n22770), .C1(conv_3[225]), .Y(n34959) );
  AOI2BB2XL U24022 ( .B0(n35195), .B1(n34962), .A0N(n34959), .A1N(n16672), .Y(
        n19267) );
  AOI22XL U24023 ( .A0(n16666), .A1(conv_3[165]), .B0(n16673), .B1(conv_3[195]), .Y(n19263) );
  NAND2XL U24024 ( .A(n19263), .B(n19262), .Y(n34955) );
  AOI22XL U24025 ( .A0(n20978), .A1(conv_3[285]), .B0(n22690), .B1(conv_3[270]), .Y(n19265) );
  NAND2XL U24026 ( .A(n19265), .B(n19264), .Y(n34960) );
  AOI22XL U24027 ( .A0(n16660), .A1(n34955), .B0(n16671), .B1(n34960), .Y(
        n19266) );
  OAI211XL U24028 ( .A0(n25853), .A1(n34968), .B0(n19267), .C0(n19266), .Y(
        n19268) );
  AOI211XL U24029 ( .A0(n16755), .A1(n34972), .B0(n19269), .C0(n19268), .Y(
        n19608) );
  NAND2XL U24030 ( .A(n26470), .B(n21831), .Y(n25872) );
  AOI22XL U24031 ( .A0(n26081), .A1(n21235), .B0(n26276), .B1(n19280), .Y(
        n19270) );
  OAI21XL U24032 ( .A0(n21236), .A1(n25987), .B0(n19270), .Y(n19292) );
  AOI22XL U24033 ( .A0(n16716), .A1(conv_3[65]), .B0(n22759), .B1(conv_3[35]), 
        .Y(n19272) );
  AOI22XL U24034 ( .A0(n16666), .A1(conv_3[50]), .B0(n18240), .B1(conv_3[80]), 
        .Y(n19271) );
  NAND2XL U24035 ( .A(n19272), .B(n19271), .Y(n21241) );
  INVXL U24036 ( .A(n34903), .Y(n26086) );
  INVXL U24037 ( .A(conv_3[305]), .Y(n31448) );
  INVXL U24038 ( .A(conv_3[275]), .Y(n31732) );
  OAI22XL U24039 ( .A0(n22612), .A1(n31448), .B0(n22717), .B1(n31732), .Y(
        n19274) );
  INVXL U24040 ( .A(conv_3[290]), .Y(n31881) );
  INVXL U24041 ( .A(conv_3[320]), .Y(n31906) );
  OAI22XL U24042 ( .A0(n22546), .A1(n31881), .B0(n18321), .B1(n31906), .Y(
        n19273) );
  OAI22XL U24043 ( .A0(n21238), .A1(n26086), .B0(n21243), .B1(n26474), .Y(
        n19275) );
  AOI21XL U24044 ( .A0(n35195), .A1(n21241), .B0(n19275), .Y(n19290) );
  AOI22XL U24045 ( .A0(n22021), .A1(conv_3[425]), .B0(n21887), .B1(conv_3[440]), .Y(n19279) );
  AOI22XL U24046 ( .A0(n16734), .A1(conv_3[410]), .B0(n21991), .B1(n20503), 
        .Y(n19278) );
  AOI22XL U24047 ( .A0(n21954), .A1(conv_3[395]), .B0(n22015), .B1(conv_3[20]), 
        .Y(n19277) );
  NAND2XL U24048 ( .A(n21992), .B(conv_3[5]), .Y(n19276) );
  NAND4XL U24049 ( .A(n19279), .B(n19278), .C(n19277), .D(n19276), .Y(n20508)
         );
  INVXL U24050 ( .A(N17708), .Y(n21688) );
  AOI2BB1XL U24051 ( .A0N(n21236), .A1N(n21688), .B0(n19280), .Y(n21246) );
  OAI22XL U24052 ( .A0(n19902), .A1(n31589), .B0(n22612), .B1(n31619), .Y(
        n19281) );
  OAI22XL U24053 ( .A0(n35143), .A1(n21246), .B0(n21244), .B1(n35198), .Y(
        n19288) );
  INVXL U24054 ( .A(conv_3[95]), .Y(n31684) );
  OAI22XL U24055 ( .A0(n16668), .A1(n31684), .B0(n24039), .B1(n34400), .Y(
        n19284) );
  INVXL U24056 ( .A(conv_3[110]), .Y(n31773) );
  OAI22XL U24057 ( .A0(n19401), .A1(n31773), .B0(n22612), .B1(n31403), .Y(
        n19283) );
  INVXL U24058 ( .A(conv_3[350]), .Y(n31484) );
  INVXL U24059 ( .A(conv_3[365]), .Y(n31641) );
  OAI22XL U24060 ( .A0(n19902), .A1(n31484), .B0(n22612), .B1(n31641), .Y(
        n19285) );
  AOI211XL U24061 ( .A0(conv_3[335]), .A1(n22616), .B0(n19286), .C0(n19285), 
        .Y(n21253) );
  OAI22XL U24062 ( .A0(n21245), .A1(n18208), .B0(n21253), .B1(n26039), .Y(
        n19287) );
  AOI211XL U24063 ( .A0(n16755), .A1(n20508), .B0(n19288), .C0(n19287), .Y(
        n19289) );
  OAI211XL U24064 ( .A0(n29160), .A1(n26085), .B0(n19290), .C0(n19289), .Y(
        n19291) );
  AOI211XL U24065 ( .A0(conv_3[215]), .A1(n26082), .B0(n19292), .C0(n19291), 
        .Y(n19600) );
  AOI22XL U24066 ( .A0(n16666), .A1(conv_3[296]), .B0(n22759), .B1(conv_3[281]), .Y(n19293) );
  NAND2XL U24067 ( .A(n19294), .B(n19293), .Y(n21306) );
  AOI22XL U24068 ( .A0(n16671), .A1(n21306), .B0(n35231), .B1(n21305), .Y(
        n19314) );
  NAND2XL U24069 ( .A(n26276), .B(n21688), .Y(n26026) );
  NAND2XL U24070 ( .A(n19296), .B(n19295), .Y(n21307) );
  AOI22XL U24071 ( .A0(n16659), .A1(n21319), .B0(n35195), .B1(n21307), .Y(
        n19300) );
  AOI22XL U24072 ( .A0(n16666), .A1(conv_3[116]), .B0(n16662), .B1(conv_3[131]), .Y(n19297) );
  NAND2XL U24073 ( .A(n19298), .B(n19297), .Y(n21320) );
  NAND2XL U24074 ( .A(n35236), .B(n21320), .Y(n19299) );
  OAI211XL U24075 ( .A0(n21313), .A1(n26026), .B0(n19300), .C0(n19299), .Y(
        n19313) );
  INVXL U24076 ( .A(conv_3[341]), .Y(n31969) );
  INVXL U24077 ( .A(conv_3[356]), .Y(n31472) );
  OAI22XL U24078 ( .A0(n19401), .A1(n31472), .B0(n22612), .B1(n31635), .Y(
        n19301) );
  AOI211XL U24079 ( .A0(conv_3[386]), .A1(n16673), .B0(n19302), .C0(n19301), 
        .Y(n21310) );
  INVXL U24080 ( .A(conv_3[206]), .Y(n31858) );
  INVXL U24081 ( .A(conv_3[191]), .Y(n31606) );
  OAI22XL U24082 ( .A0(n22612), .A1(n31606), .B0(n22717), .B1(n32320), .Y(
        n19303) );
  AOI211XL U24083 ( .A0(conv_3[176]), .A1(n21011), .B0(n19304), .C0(n19303), 
        .Y(n21317) );
  OAI22XL U24084 ( .A0(n21310), .A1(n26039), .B0(n21317), .B1(n35198), .Y(
        n19312) );
  INVXL U24085 ( .A(conv_3[431]), .Y(n31730) );
  OAI22XL U24086 ( .A0(n19416), .A1(n31730), .B0(n16669), .B1(n32042), .Y(
        n19308) );
  AOI22XL U24087 ( .A0(n16734), .A1(conv_3[416]), .B0(n21991), .B1(n21314), 
        .Y(n19306) );
  AOI22XL U24088 ( .A0(n21887), .A1(conv_3[446]), .B0(conv_3[26]), .B1(n22015), 
        .Y(n19305) );
  NAND2XL U24089 ( .A(n19306), .B(n19305), .Y(n19307) );
  AOI211XL U24090 ( .A0(n21992), .A1(conv_3[11]), .B0(n19308), .C0(n19307), 
        .Y(n20577) );
  AOI22XL U24091 ( .A0(conv_3[236]), .A1(n26059), .B0(n34903), .B1(n21314), 
        .Y(n19310) );
  AOI22XL U24092 ( .A0(conv_3[221]), .A1(n26082), .B0(n26081), .B1(n21318), 
        .Y(n19309) );
  OAI211XL U24093 ( .A0(n20577), .A1(n35159), .B0(n19310), .C0(n19309), .Y(
        n19311) );
  NOR4BXL U24094 ( .AN(n19314), .B(n19313), .C(n19312), .D(n19311), .Y(n19597)
         );
  AOI22XL U24095 ( .A0(n22021), .A1(conv_3[426]), .B0(n21887), .B1(conv_3[441]), .Y(n19318) );
  AOI22XL U24096 ( .A0(n16734), .A1(conv_3[411]), .B0(n21991), .B1(n21270), 
        .Y(n19317) );
  AOI22XL U24097 ( .A0(n21954), .A1(conv_3[396]), .B0(conv_3[21]), .B1(n22015), 
        .Y(n19316) );
  NAND2XL U24098 ( .A(n21992), .B(conv_3[6]), .Y(n19315) );
  NAND4XL U24099 ( .A(n19318), .B(n19317), .C(n19316), .D(n19315), .Y(n20462)
         );
  INVXL U24100 ( .A(conv_3[231]), .Y(n32093) );
  AOI22XL U24101 ( .A0(n16666), .A1(conv_3[111]), .B0(n18658), .B1(conv_3[96]), 
        .Y(n19319) );
  NAND2XL U24102 ( .A(n19320), .B(n19319), .Y(n21258) );
  AOI22XL U24103 ( .A0(n35236), .A1(n21258), .B0(n26081), .B1(n21265), .Y(
        n19321) );
  OAI21XL U24104 ( .A0(n32093), .A1(n26085), .B0(n19321), .Y(n19335) );
  INVXL U24105 ( .A(n26026), .Y(n25875) );
  AOI22XL U24106 ( .A0(n34903), .A1(n21270), .B0(n25875), .B1(n21263), .Y(
        n19333) );
  AOI22XL U24107 ( .A0(n16666), .A1(conv_3[351]), .B0(n16662), .B1(conv_3[366]), .Y(n19323) );
  NAND2XL U24108 ( .A(n19323), .B(n19322), .Y(n21259) );
  AOI22XL U24109 ( .A0(conv_3[216]), .A1(n26082), .B0(n19179), .B1(n21259), 
        .Y(n19332) );
  AOI22XL U24110 ( .A0(n16666), .A1(conv_3[51]), .B0(n16662), .B1(conv_3[66]), 
        .Y(n19325) );
  NAND2XL U24111 ( .A(n19325), .B(n19324), .Y(n21271) );
  NAND2XL U24112 ( .A(n35143), .B(n25987), .Y(n25879) );
  INVXL U24113 ( .A(n25879), .Y(n25975) );
  AOI2BB2XL U24114 ( .B0(n35195), .B1(n21271), .A0N(n25975), .A1N(n21262), .Y(
        n19331) );
  AOI22XL U24115 ( .A0(n16662), .A1(conv_3[186]), .B0(n18240), .B1(conv_3[201]), .Y(n19327) );
  AOI22XL U24116 ( .A0(n16666), .A1(conv_3[171]), .B0(n25299), .B1(conv_3[156]), .Y(n19326) );
  NAND2XL U24117 ( .A(n19327), .B(n19326), .Y(n21266) );
  AOI22XL U24118 ( .A0(n16666), .A1(conv_3[291]), .B0(n16662), .B1(conv_3[306]), .Y(n19329) );
  NAND2XL U24119 ( .A(n19329), .B(n19328), .Y(n21257) );
  AOI22XL U24120 ( .A0(n16660), .A1(n21266), .B0(n16671), .B1(n21257), .Y(
        n19330) );
  NAND4XL U24121 ( .A(n19333), .B(n19332), .C(n19331), .D(n19330), .Y(n19334)
         );
  AOI211XL U24122 ( .A0(n16755), .A1(n20462), .B0(n19335), .C0(n19334), .Y(
        n19596) );
  NAND2XL U24123 ( .A(n19337), .B(n19336), .Y(n21288) );
  AOI22XL U24124 ( .A0(n16666), .A1(conv_3[294]), .B0(n16662), .B1(conv_3[309]), .Y(n19339) );
  NAND2XL U24125 ( .A(n19339), .B(n19338), .Y(n21287) );
  AOI22XL U24126 ( .A0(n16660), .A1(n21288), .B0(n16671), .B1(n21287), .Y(
        n19357) );
  INVXL U24127 ( .A(conv_3[354]), .Y(n31490) );
  OAI22XL U24128 ( .A0(n19902), .A1(n31490), .B0(n18321), .B1(n31506), .Y(
        n19341) );
  INVXL U24129 ( .A(conv_3[339]), .Y(n31957) );
  OAI22XL U24130 ( .A0(n22612), .A1(n35763), .B0(n22717), .B1(n31957), .Y(
        n19340) );
  AOI22XL U24131 ( .A0(conv_3[234]), .A1(n26059), .B0(conv_3[219]), .B1(n26082), .Y(n19345) );
  AOI22XL U24132 ( .A0(n16666), .A1(conv_3[114]), .B0(n16662), .B1(conv_3[129]), .Y(n19343) );
  AOI22XL U24133 ( .A0(n22759), .A1(conv_3[99]), .B0(n16673), .B1(conv_3[144]), 
        .Y(n19342) );
  NAND2XL U24134 ( .A(n19343), .B(n19342), .Y(n21304) );
  NAND2XL U24135 ( .A(n35236), .B(n21304), .Y(n19344) );
  OAI211XL U24136 ( .A0(n21285), .A1(n26039), .B0(n19345), .C0(n19344), .Y(
        n19356) );
  INVXL U24137 ( .A(conv_3[54]), .Y(n31198) );
  INVXL U24138 ( .A(conv_3[69]), .Y(n31478) );
  OAI22XL U24139 ( .A0(n22546), .A1(n31198), .B0(n22612), .B1(n31478), .Y(
        n19347) );
  INVXL U24140 ( .A(conv_3[39]), .Y(n31231) );
  INVXL U24141 ( .A(conv_3[84]), .Y(n35609) );
  OAI22XL U24142 ( .A0(n22717), .A1(n31231), .B0(n18321), .B1(n35609), .Y(
        n19346) );
  OAI22XL U24143 ( .A0(n35143), .A1(n21289), .B0(n21290), .B1(n35239), .Y(
        n19355) );
  INVXL U24144 ( .A(conv_3[444]), .Y(n35791) );
  OAI22XL U24145 ( .A0(n21810), .A1(n35791), .B0(n16669), .B1(n32047), .Y(
        n19351) );
  AOI22XL U24146 ( .A0(n22021), .A1(conv_3[429]), .B0(n21991), .B1(n21282), 
        .Y(n19349) );
  AOI22XL U24147 ( .A0(n16734), .A1(conv_3[414]), .B0(conv_3[24]), .B1(n22015), 
        .Y(n19348) );
  NAND2XL U24148 ( .A(n19349), .B(n19348), .Y(n19350) );
  AOI211XL U24149 ( .A0(n21992), .A1(conv_3[9]), .B0(n19351), .C0(n19350), .Y(
        n20578) );
  AOI22XL U24150 ( .A0(n26081), .A1(n21297), .B0(n34903), .B1(n21282), .Y(
        n19353) );
  AOI22XL U24151 ( .A0(n26066), .A1(n21286), .B0(n25875), .B1(n21295), .Y(
        n19352) );
  OAI211XL U24152 ( .A0(n20578), .A1(n35159), .B0(n19353), .C0(n19352), .Y(
        n19354) );
  NOR4BXL U24153 ( .AN(n19357), .B(n19356), .C(n19355), .D(n19354), .Y(n19595)
         );
  NAND4XL U24154 ( .A(n19600), .B(n19597), .C(n19596), .D(n19595), .Y(n19522)
         );
  INVXL U24155 ( .A(pool[129]), .Y(n19742) );
  AOI22XL U24156 ( .A0(n21887), .A1(conv_3[439]), .B0(n21991), .B1(n21201), 
        .Y(n19361) );
  AOI22XL U24157 ( .A0(n16734), .A1(conv_3[409]), .B0(n21954), .B1(conv_3[394]), .Y(n19360) );
  AOI22XL U24158 ( .A0(n22021), .A1(conv_3[424]), .B0(n22015), .B1(conv_3[19]), 
        .Y(n19359) );
  NAND2XL U24159 ( .A(n21992), .B(conv_3[4]), .Y(n19358) );
  NAND4XL U24160 ( .A(n19361), .B(n19360), .C(n19359), .D(n19358), .Y(n20498)
         );
  INVXL U24161 ( .A(conv_3[34]), .Y(n29668) );
  INVXL U24162 ( .A(conv_3[49]), .Y(n23211) );
  OAI22XL U24163 ( .A0(n22546), .A1(n23211), .B0(n22612), .B1(n23904), .Y(
        n19362) );
  AOI211XL U24164 ( .A0(conv_3[79]), .A1(n18240), .B0(n19363), .C0(n19362), 
        .Y(n21192) );
  AOI22XL U24165 ( .A0(n16716), .A1(conv_3[304]), .B0(n16673), .B1(conv_3[319]), .Y(n19365) );
  AOI22XL U24166 ( .A0(n16666), .A1(conv_3[289]), .B0(n22690), .B1(conv_3[274]), .Y(n19364) );
  NAND2XL U24167 ( .A(n19365), .B(n19364), .Y(n21190) );
  AOI22XL U24168 ( .A0(n16671), .A1(n21190), .B0(n34903), .B1(n21201), .Y(
        n19369) );
  AOI22XL U24169 ( .A0(n16666), .A1(conv_3[109]), .B0(n18658), .B1(conv_3[94]), 
        .Y(n19367) );
  NAND2XL U24170 ( .A(n19367), .B(n19366), .Y(n21196) );
  NAND2XL U24171 ( .A(n35236), .B(n21196), .Y(n19368) );
  OAI211XL U24172 ( .A0(n21192), .A1(n35239), .B0(n19369), .C0(n19368), .Y(
        n19379) );
  INVXL U24173 ( .A(n20490), .Y(n21194) );
  AOI22XL U24174 ( .A0(n26081), .A1(n21195), .B0(n26066), .B1(n21194), .Y(
        n19377) );
  AOI22XL U24175 ( .A0(conv_3[229]), .A1(n26059), .B0(conv_3[214]), .B1(n26082), .Y(n19376) );
  AOI22XL U24176 ( .A0(n16666), .A1(conv_3[169]), .B0(n25299), .B1(conv_3[154]), .Y(n19370) );
  NAND2XL U24177 ( .A(n19371), .B(n19370), .Y(n21197) );
  INVXL U24178 ( .A(n21195), .Y(n20492) );
  AOI22XL U24179 ( .A0(n16660), .A1(n21197), .B0(n26276), .B1(n21191), .Y(
        n19375) );
  AOI22XL U24180 ( .A0(n16716), .A1(conv_3[364]), .B0(n22690), .B1(conv_3[334]), .Y(n19373) );
  AOI22XL U24181 ( .A0(n16666), .A1(conv_3[349]), .B0(n18240), .B1(conv_3[379]), .Y(n19372) );
  AND2XL U24182 ( .A(n19373), .B(n19372), .Y(n21193) );
  AOI2BB2XL U24183 ( .B0(n21202), .B1(n35231), .A0N(n21193), .A1N(n26039), .Y(
        n19374) );
  NAND4XL U24184 ( .A(n19377), .B(n19376), .C(n19375), .D(n19374), .Y(n19378)
         );
  AOI211XL U24185 ( .A0(n16755), .A1(n20498), .B0(n19379), .C0(n19378), .Y(
        n19741) );
  AOI22XL U24186 ( .A0(n16734), .A1(conv_3[412]), .B0(n21991), .B1(n21217), 
        .Y(n19383) );
  AOI22XL U24187 ( .A0(n22021), .A1(conv_3[427]), .B0(n21954), .B1(conv_3[397]), .Y(n19382) );
  AOI22XL U24188 ( .A0(n21887), .A1(conv_3[442]), .B0(n21992), .B1(conv_3[7]), 
        .Y(n19381) );
  NAND2XL U24189 ( .A(conv_3[22]), .B(n22015), .Y(n19380) );
  NAND4XL U24190 ( .A(n19383), .B(n19382), .C(n19381), .D(n19380), .Y(n20471)
         );
  AOI22XL U24191 ( .A0(conv_3[217]), .A1(n26082), .B0(n26081), .B1(n21228), 
        .Y(n19384) );
  OAI21XL U24192 ( .A0(n25975), .A1(n21216), .B0(n19384), .Y(n19400) );
  AOI22XL U24193 ( .A0(n34903), .A1(n21217), .B0(n25875), .B1(n21226), .Y(
        n19398) );
  AOI22XL U24194 ( .A0(n16666), .A1(conv_3[52]), .B0(n22759), .B1(conv_3[37]), 
        .Y(n19386) );
  NAND2XL U24195 ( .A(n19386), .B(n19385), .Y(n21229) );
  AOI22XL U24196 ( .A0(n35195), .A1(n21229), .B0(conv_3[232]), .B1(n26059), 
        .Y(n19397) );
  AOI22XL U24197 ( .A0(n16666), .A1(conv_3[112]), .B0(n18240), .B1(conv_3[142]), .Y(n19388) );
  AOI22XL U24198 ( .A0(n16662), .A1(conv_3[127]), .B0(n22690), .B1(conv_3[97]), 
        .Y(n19387) );
  NAND2XL U24199 ( .A(n19388), .B(n19387), .Y(n21218) );
  AOI22XL U24200 ( .A0(n16662), .A1(conv_3[307]), .B0(n22690), .B1(conv_3[277]), .Y(n19390) );
  AOI22XL U24201 ( .A0(n16666), .A1(conv_3[292]), .B0(n18240), .B1(conv_3[322]), .Y(n19389) );
  NAND2XL U24202 ( .A(n19390), .B(n19389), .Y(n21212) );
  AOI22XL U24203 ( .A0(n35236), .A1(n21218), .B0(n16671), .B1(n21212), .Y(
        n19396) );
  AOI22XL U24204 ( .A0(n16666), .A1(conv_3[172]), .B0(n16673), .B1(conv_3[202]), .Y(n19392) );
  AOI22XL U24205 ( .A0(n16662), .A1(conv_3[187]), .B0(n22759), .B1(conv_3[157]), .Y(n19391) );
  NAND2XL U24206 ( .A(n19392), .B(n19391), .Y(n21225) );
  AOI22XL U24207 ( .A0(n16662), .A1(conv_3[367]), .B0(n22690), .B1(conv_3[337]), .Y(n19393) );
  NAND2XL U24208 ( .A(n19394), .B(n19393), .Y(n21211) );
  AOI22XL U24209 ( .A0(n16660), .A1(n21225), .B0(n19179), .B1(n21211), .Y(
        n19395) );
  NAND4XL U24210 ( .A(n19398), .B(n19397), .C(n19396), .D(n19395), .Y(n19399)
         );
  AOI211XL U24211 ( .A0(n16755), .A1(n20471), .B0(n19400), .C0(n19399), .Y(
        n19591) );
  INVXL U24212 ( .A(conv_3[293]), .Y(n35722) );
  INVXL U24213 ( .A(conv_3[278]), .Y(n31743) );
  INVXL U24214 ( .A(conv_3[323]), .Y(n35742) );
  OAI22XL U24215 ( .A0(n22550), .A1(n31743), .B0(n18321), .B1(n35742), .Y(
        n19402) );
  OAI22XL U24216 ( .A0(n35143), .A1(n21343), .B0(n21339), .B1(n26474), .Y(
        n19415) );
  AOI22XL U24217 ( .A0(n28528), .A1(n21329), .B0(conv_3[233]), .B1(n26059), 
        .Y(n19414) );
  AOI22XL U24218 ( .A0(n16716), .A1(conv_3[68]), .B0(n18240), .B1(conv_3[83]), 
        .Y(n19405) );
  AOI22XL U24219 ( .A0(n16666), .A1(conv_3[53]), .B0(n25299), .B1(conv_3[38]), 
        .Y(n19404) );
  NAND2XL U24220 ( .A(n19405), .B(n19404), .Y(n21346) );
  AOI22XL U24221 ( .A0(n16666), .A1(conv_3[173]), .B0(n16662), .B1(conv_3[188]), .Y(n19407) );
  NAND2XL U24222 ( .A(n19407), .B(n19406), .Y(n21335) );
  AOI22XL U24223 ( .A0(n35195), .A1(n21346), .B0(n16660), .B1(n21335), .Y(
        n19413) );
  AOI22XL U24224 ( .A0(n16666), .A1(conv_3[113]), .B0(n16662), .B1(conv_3[128]), .Y(n19409) );
  NAND2XL U24225 ( .A(n19409), .B(n19408), .Y(n21336) );
  AOI22XL U24226 ( .A0(n16716), .A1(conv_3[368]), .B0(n22616), .B1(conv_3[338]), .Y(n19410) );
  NAND2XL U24227 ( .A(n19411), .B(n19410), .Y(n21334) );
  AOI22XL U24228 ( .A0(n35236), .A1(n21336), .B0(n19179), .B1(n21334), .Y(
        n19412) );
  NAND4BXL U24229 ( .AN(n19415), .B(n19414), .C(n19413), .D(n19412), .Y(n19424) );
  INVXL U24230 ( .A(conv_3[428]), .Y(n31706) );
  INVXL U24231 ( .A(conv_3[443]), .Y(n32112) );
  OAI22XL U24232 ( .A0(n19416), .A1(n31706), .B0(n21810), .B1(n32112), .Y(
        n19420) );
  AOI22XL U24233 ( .A0(n21954), .A1(conv_3[398]), .B0(n21991), .B1(n21340), 
        .Y(n19418) );
  AOI22XL U24234 ( .A0(n16734), .A1(conv_3[413]), .B0(conv_3[23]), .B1(n22015), 
        .Y(n19417) );
  NAND2XL U24235 ( .A(n19418), .B(n19417), .Y(n19419) );
  AOI211XL U24236 ( .A0(n21992), .A1(conv_3[8]), .B0(n19420), .C0(n19419), .Y(
        n20581) );
  AOI22XL U24237 ( .A0(n26081), .A1(n21333), .B0(n26276), .B1(n21331), .Y(
        n19422) );
  AOI22XL U24238 ( .A0(conv_3[218]), .A1(n26082), .B0(n34903), .B1(n21340), 
        .Y(n19421) );
  OAI211XL U24239 ( .A0(n20581), .A1(n35159), .B0(n19422), .C0(n19421), .Y(
        n19423) );
  INVXL U24240 ( .A(conv_3[145]), .Y(n33469) );
  INVXL U24241 ( .A(conv_3[130]), .Y(n33799) );
  OAI22XL U24242 ( .A0(n22740), .A1(n33799), .B0(n22717), .B1(n31672), .Y(
        n19425) );
  OAI22XL U24243 ( .A0(n19427), .A1(n25872), .B0(n21356), .B1(n18208), .Y(
        n19447) );
  INVXL U24244 ( .A(conv_3[370]), .Y(n33835) );
  INVXL U24245 ( .A(conv_3[355]), .Y(n33476) );
  INVXL U24246 ( .A(conv_3[385]), .Y(n31465) );
  OAI22XL U24247 ( .A0(n19902), .A1(n33476), .B0(n18321), .B1(n31465), .Y(
        n19428) );
  AOI211XL U24248 ( .A0(conv_3[340]), .A1(n22759), .B0(n19429), .C0(n19428), 
        .Y(n21352) );
  NAND2XL U24249 ( .A(n19431), .B(n19430), .Y(n21364) );
  AOI22XL U24250 ( .A0(n22759), .A1(conv_3[280]), .B0(n18240), .B1(conv_3[325]), .Y(n19433) );
  NAND2XL U24251 ( .A(n19433), .B(n19432), .Y(n21361) );
  AOI22XL U24252 ( .A0(n16660), .A1(n21364), .B0(n16671), .B1(n21361), .Y(
        n19435) );
  NAND2XL U24253 ( .A(n25879), .B(n21363), .Y(n19434) );
  OAI211XL U24254 ( .A0(n21352), .A1(n26039), .B0(n19435), .C0(n19434), .Y(
        n19446) );
  OAI22XL U24255 ( .A0(n19436), .A1(n22014), .B0(n31256), .B1(n21953), .Y(
        n19440) );
  AOI22XL U24256 ( .A0(n16734), .A1(conv_3[415]), .B0(n21887), .B1(conv_3[445]), .Y(n19438) );
  AOI22XL U24257 ( .A0(n22021), .A1(conv_3[430]), .B0(n21954), .B1(conv_3[400]), .Y(n19437) );
  NAND2XL U24258 ( .A(n19438), .B(n19437), .Y(n19439) );
  AOI211XL U24259 ( .A0(n21992), .A1(conv_3[10]), .B0(n19440), .C0(n19439), 
        .Y(n20588) );
  AOI22XL U24260 ( .A0(conv_3[220]), .A1(n26082), .B0(n26276), .B1(n20481), 
        .Y(n19444) );
  AOI22XL U24261 ( .A0(n16662), .A1(conv_3[70]), .B0(n22690), .B1(conv_3[40]), 
        .Y(n19441) );
  NAND2XL U24262 ( .A(n19442), .B(n19441), .Y(n21362) );
  AOI22XL U24263 ( .A0(n35195), .A1(n21362), .B0(n34903), .B1(n21353), .Y(
        n19443) );
  OAI211XL U24264 ( .A0(n20588), .A1(n35159), .B0(n19444), .C0(n19443), .Y(
        n19445) );
  NOR4XL U24265 ( .A(n19448), .B(n19447), .C(n19446), .D(n19445), .Y(n19601)
         );
  NAND4XL U24266 ( .A(n19741), .B(n19591), .C(n19590), .D(n19601), .Y(n19521)
         );
  AOI22XL U24267 ( .A0(n21990), .A1(conv_3[423]), .B0(n21954), .B1(conv_3[393]), .Y(n19452) );
  AOI22XL U24268 ( .A0(n16734), .A1(conv_3[408]), .B0(n21887), .B1(conv_3[438]), .Y(n19451) );
  AOI22XL U24269 ( .A0(n21991), .A1(n21124), .B0(n22015), .B1(conv_3[18]), .Y(
        n19450) );
  NAND2XL U24270 ( .A(n21992), .B(conv_3[3]), .Y(n19449) );
  NAND4XL U24271 ( .A(n19452), .B(n19451), .C(n19450), .D(n19449), .Y(n20429)
         );
  INVXL U24272 ( .A(conv_3[228]), .Y(n29674) );
  AOI22XL U24273 ( .A0(n16666), .A1(conv_3[108]), .B0(n16673), .B1(conv_3[138]), .Y(n19453) );
  NAND2XL U24274 ( .A(n19454), .B(n19453), .Y(n21135) );
  AOI22XL U24275 ( .A0(n35236), .A1(n21135), .B0(n26081), .B1(n21130), .Y(
        n19455) );
  OAI21XL U24276 ( .A0(n29674), .A1(n26085), .B0(n19455), .Y(n19469) );
  AOI22XL U24277 ( .A0(n34903), .A1(n21124), .B0(n21132), .B1(n25879), .Y(
        n19467) );
  AOI2BB2XL U24278 ( .B0(n20422), .B1(n22713), .A0N(n21688), .A1N(n21130), .Y(
        n21131) );
  AOI22XL U24279 ( .A0(n26082), .A1(conv_3[213]), .B0(n26276), .B1(n21131), 
        .Y(n19466) );
  AOI22XL U24280 ( .A0(n16666), .A1(conv_3[48]), .B0(n22690), .B1(conv_3[33]), 
        .Y(n19456) );
  NAND2XL U24281 ( .A(n19457), .B(n19456), .Y(n21134) );
  AOI22XL U24282 ( .A0(n16666), .A1(conv_3[348]), .B0(n22690), .B1(conv_3[333]), .Y(n19458) );
  NAND2XL U24283 ( .A(n19459), .B(n19458), .Y(n21125) );
  AOI22XL U24284 ( .A0(n35195), .A1(n21134), .B0(n19179), .B1(n21125), .Y(
        n19465) );
  AOI22XL U24285 ( .A0(n16666), .A1(conv_3[168]), .B0(n22759), .B1(conv_3[153]), .Y(n19461) );
  AOI22XL U24286 ( .A0(n16662), .A1(conv_3[183]), .B0(n16673), .B1(conv_3[198]), .Y(n19460) );
  NAND2XL U24287 ( .A(n19461), .B(n19460), .Y(n21126) );
  AOI22XL U24288 ( .A0(n16666), .A1(conv_3[288]), .B0(n22690), .B1(conv_3[273]), .Y(n19463) );
  NAND2XL U24289 ( .A(n19463), .B(n19462), .Y(n21133) );
  AOI22XL U24290 ( .A0(n16660), .A1(n21126), .B0(n16671), .B1(n21133), .Y(
        n19464) );
  NAND4XL U24291 ( .A(n19467), .B(n19466), .C(n19465), .D(n19464), .Y(n19468)
         );
  INVXL U24292 ( .A(pool[127]), .Y(n35025) );
  AOI211XL U24293 ( .A0(n21167), .A1(n28292), .B0(n21173), .C0(n19474), .Y(
        n20441) );
  NAND2XL U24294 ( .A(n19473), .B(n19472), .Y(n21177) );
  INVXL U24295 ( .A(conv_3[227]), .Y(n30850) );
  OAI21XL U24296 ( .A0(n21167), .A1(n20433), .B0(n28528), .Y(n19477) );
  AOI32XL U24297 ( .A0(conv_3[212]), .A1(n23055), .A2(n19475), .B0(n19474), 
        .B1(n23055), .Y(n19476) );
  OAI211XL U24298 ( .A0(n26085), .A1(n30850), .B0(n19477), .C0(n19476), .Y(
        n19491) );
  INVXL U24299 ( .A(conv_3[407]), .Y(n30548) );
  OAI22XL U24300 ( .A0(n21172), .A1(n22014), .B0(n21944), .B1(n30548), .Y(
        n19481) );
  AOI22XL U24301 ( .A0(n21887), .A1(conv_3[437]), .B0(n21954), .B1(conv_3[392]), .Y(n19479) );
  AOI22XL U24302 ( .A0(n22021), .A1(conv_3[422]), .B0(n22015), .B1(conv_3[17]), 
        .Y(n19478) );
  NAND2XL U24303 ( .A(n19479), .B(n19478), .Y(n19480) );
  AOI211XL U24304 ( .A0(n21992), .A1(conv_3[2]), .B0(n19481), .C0(n19480), .Y(
        n20436) );
  OR2XL U24305 ( .A(n21173), .B(n21167), .Y(n21170) );
  AOI22XL U24306 ( .A0(n16666), .A1(conv_3[347]), .B0(n16662), .B1(conv_3[362]), .Y(n19482) );
  NAND2XL U24307 ( .A(n19483), .B(n19482), .Y(n21168) );
  AOI22XL U24308 ( .A0(n34906), .A1(n21170), .B0(n19179), .B1(n21168), .Y(
        n19489) );
  AOI22XL U24309 ( .A0(n20978), .A1(conv_3[107]), .B0(n16662), .B1(conv_3[122]), .Y(n19485) );
  NAND2XL U24310 ( .A(n19485), .B(n19484), .Y(n21175) );
  AOI22XL U24311 ( .A0(n22690), .A1(conv_3[152]), .B0(n16673), .B1(conv_3[197]), .Y(n19487) );
  AOI22XL U24312 ( .A0(n20978), .A1(conv_3[167]), .B0(n16662), .B1(conv_3[182]), .Y(n19486) );
  NAND2XL U24313 ( .A(n19487), .B(n19486), .Y(n21169) );
  AOI22XL U24314 ( .A0(n35236), .A1(n21175), .B0(n16660), .B1(n21169), .Y(
        n19488) );
  OAI211XL U24315 ( .A0(n20436), .A1(n35159), .B0(n19489), .C0(n19488), .Y(
        n19490) );
  AOI211XL U24316 ( .A0(n35195), .A1(n21177), .B0(n19491), .C0(n19490), .Y(
        n19495) );
  AOI22XL U24317 ( .A0(n16666), .A1(conv_3[287]), .B0(n16662), .B1(conv_3[302]), .Y(n19492) );
  NAND2XL U24318 ( .A(n19493), .B(n19492), .Y(n21176) );
  NAND2XL U24319 ( .A(n16671), .B(n21176), .Y(n19494) );
  AOI22XL U24320 ( .A0(n22021), .A1(conv_3[421]), .B0(n16734), .B1(conv_3[406]), .Y(n19499) );
  AOI22XL U24321 ( .A0(n21887), .A1(conv_3[436]), .B0(n21991), .B1(n21144), 
        .Y(n19498) );
  AOI22XL U24322 ( .A0(n21954), .A1(conv_3[391]), .B0(n22015), .B1(conv_3[16]), 
        .Y(n19497) );
  NAND2XL U24323 ( .A(n21992), .B(conv_3[1]), .Y(n19496) );
  NAND4XL U24324 ( .A(n19499), .B(n19498), .C(n19497), .D(n19496), .Y(n20451)
         );
  AOI22XL U24325 ( .A0(conv_3[226]), .A1(n26059), .B0(n26081), .B1(n21150), 
        .Y(n19501) );
  NAND2XL U24326 ( .A(n26082), .B(conv_3[211]), .Y(n19500) );
  OAI211XL U24327 ( .A0(n21147), .A1(n26026), .B0(n19501), .C0(n19500), .Y(
        n19517) );
  AOI2BB2XL U24328 ( .B0(n34903), .B1(n21144), .A0N(n25987), .A1N(n21148), .Y(
        n19515) );
  AOI22XL U24329 ( .A0(n20978), .A1(conv_3[106]), .B0(n22690), .B1(conv_3[91]), 
        .Y(n19502) );
  NAND2XL U24330 ( .A(n19503), .B(n19502), .Y(n21151) );
  AOI22XL U24331 ( .A0(n35236), .A1(n21151), .B0(n35231), .B1(n21155), .Y(
        n19514) );
  AOI22XL U24332 ( .A0(n16666), .A1(conv_3[166]), .B0(n22690), .B1(conv_3[151]), .Y(n19505) );
  NAND2XL U24333 ( .A(n19505), .B(n19504), .Y(n21154) );
  AOI22XL U24334 ( .A0(n16662), .A1(conv_3[361]), .B0(n22690), .B1(conv_3[331]), .Y(n19506) );
  NAND2XL U24335 ( .A(n19507), .B(n19506), .Y(n21156) );
  AOI22XL U24336 ( .A0(n16660), .A1(n21154), .B0(n19179), .B1(n21156), .Y(
        n19513) );
  AOI22XL U24337 ( .A0(n16666), .A1(conv_3[46]), .B0(n16662), .B1(conv_3[61]), 
        .Y(n19509) );
  AOI22XL U24338 ( .A0(n16662), .A1(conv_3[301]), .B0(n22690), .B1(conv_3[271]), .Y(n19511) );
  NAND2XL U24339 ( .A(n19511), .B(n19510), .Y(n21157) );
  AOI22XL U24340 ( .A0(n35195), .A1(n21158), .B0(n16671), .B1(n21157), .Y(
        n19512) );
  NAND4XL U24341 ( .A(n19515), .B(n19514), .C(n19513), .D(n19512), .Y(n19516)
         );
  AOI222XL U24342 ( .A0(pool[125]), .A1(pool[126]), .B0(pool[125]), .B1(n35023), .C0(pool[126]), .C1(n35023), .Y(n19518) );
  AOI222XL U24343 ( .A0(n35025), .A1(n35024), .B0(n35025), .B1(n19518), .C0(
        n35024), .C1(n19518), .Y(n19519) );
  AOI222XL U24344 ( .A0(n35028), .A1(pool[128]), .B0(n35028), .B1(n19519), 
        .C0(pool[128]), .C1(n19519), .Y(n19520) );
  AOI221XL U24345 ( .A0(n19522), .A1(n19742), .B0(n19521), .B1(n19742), .C0(
        n19520), .Y(n19605) );
  OAI22XL U24346 ( .A0(n22717), .A1(n32219), .B0(n22716), .B1(n32204), .Y(
        n19524) );
  INVXL U24347 ( .A(conv_3[374]), .Y(n32127) );
  OAI22XL U24348 ( .A0(n19401), .A1(n32135), .B0(n22612), .B1(n32127), .Y(
        n19523) );
  OAI22XL U24349 ( .A0(n35143), .A1(n21385), .B0(n21393), .B1(n26039), .Y(
        n19544) );
  INVXL U24350 ( .A(conv_3[209]), .Y(n32277) );
  OAI22XL U24351 ( .A0(n18286), .A1(n32226), .B0(n22716), .B1(n32277), .Y(
        n19525) );
  INVXL U24352 ( .A(conv_3[119]), .Y(n32270) );
  INVXL U24353 ( .A(conv_3[104]), .Y(n32120) );
  OAI22XL U24354 ( .A0(n19401), .A1(n32270), .B0(n22717), .B1(n32120), .Y(
        n19527) );
  OAI2BB2XL U24355 ( .B0(n21389), .B1(n18208), .A0N(n21381), .A1N(n34903), .Y(
        n19529) );
  AOI211XL U24356 ( .A0(n20542), .A1(n26276), .B0(n19530), .C0(n19529), .Y(
        n19543) );
  AOI22XL U24357 ( .A0(n16666), .A1(conv_3[59]), .B0(n16716), .B1(conv_3[74]), 
        .Y(n19532) );
  AOI22XL U24358 ( .A0(n22759), .A1(conv_3[44]), .B0(n18240), .B1(conv_3[89]), 
        .Y(n19531) );
  NAND2XL U24359 ( .A(n19532), .B(n19531), .Y(n21392) );
  NAND2XL U24360 ( .A(n19534), .B(n19533), .Y(n21387) );
  AOI22XL U24361 ( .A0(n35195), .A1(n21392), .B0(n16671), .B1(n21387), .Y(
        n19542) );
  AOI22XL U24362 ( .A0(n21887), .A1(conv_3[449]), .B0(n21991), .B1(n21381), 
        .Y(n19538) );
  AOI22XL U24363 ( .A0(n22021), .A1(conv_3[434]), .B0(n21954), .B1(conv_3[404]), .Y(n19537) );
  AOI22XL U24364 ( .A0(n16734), .A1(conv_3[419]), .B0(n21992), .B1(conv_3[14]), 
        .Y(n19536) );
  NAND2XL U24365 ( .A(conv_3[29]), .B(n22015), .Y(n19535) );
  NAND4XL U24366 ( .A(n19538), .B(n19537), .C(n19536), .D(n19535), .Y(n20545)
         );
  INVXL U24367 ( .A(conv_3[239]), .Y(n33904) );
  OAI22XL U24368 ( .A0(n20538), .A1(n25987), .B0(n33904), .B1(n26085), .Y(
        n19540) );
  INVXL U24369 ( .A(n20541), .Y(n21391) );
  INVXL U24370 ( .A(conv_3[224]), .Y(n32142) );
  OAI22XL U24371 ( .A0(n21391), .A1(n25872), .B0(n32142), .B1(n26029), .Y(
        n19539) );
  AOI211XL U24372 ( .A0(n16755), .A1(n20545), .B0(n19540), .C0(n19539), .Y(
        n19541) );
  NAND4BXL U24373 ( .AN(n19544), .B(n19543), .C(n19542), .D(n19541), .Y(n19604) );
  INVXL U24374 ( .A(conv_3[147]), .Y(n32793) );
  INVXL U24375 ( .A(conv_3[117]), .Y(n34201) );
  INVXL U24376 ( .A(conv_3[102]), .Y(n34192) );
  OAI22XL U24377 ( .A0(n19401), .A1(n34201), .B0(n16668), .B1(n34192), .Y(
        n19545) );
  INVXL U24378 ( .A(conv_3[222]), .Y(n34653) );
  OAI22XL U24379 ( .A0(n21428), .A1(n18208), .B0(n34653), .B1(n26029), .Y(
        n19547) );
  AOI21XL U24380 ( .A0(n26081), .A1(n21431), .B0(n19547), .Y(n19566) );
  INVXL U24381 ( .A(n19558), .Y(n21424) );
  AOI22XL U24382 ( .A0(n34903), .A1(n21423), .B0(n25875), .B1(n21424), .Y(
        n19565) );
  AOI22XL U24383 ( .A0(n22616), .A1(conv_3[42]), .B0(n16673), .B1(conv_3[87]), 
        .Y(n19548) );
  NAND2XL U24384 ( .A(n19549), .B(n19548), .Y(n21432) );
  AOI22XL U24385 ( .A0(n35195), .A1(n21432), .B0(conv_3[237]), .B1(n26059), 
        .Y(n19564) );
  AOI22XL U24386 ( .A0(n22021), .A1(conv_3[432]), .B0(n21887), .B1(conv_3[447]), .Y(n19553) );
  AOI22XL U24387 ( .A0(n16734), .A1(conv_3[417]), .B0(n21991), .B1(n21423), 
        .Y(n19552) );
  AOI22XL U24388 ( .A0(n21954), .A1(conv_3[402]), .B0(conv_3[27]), .B1(n22015), 
        .Y(n19551) );
  NAND2XL U24389 ( .A(n21992), .B(conv_3[12]), .Y(n19550) );
  NAND4XL U24390 ( .A(n19553), .B(n19552), .C(n19551), .D(n19550), .Y(n20568)
         );
  INVXL U24391 ( .A(conv_3[312]), .Y(n33110) );
  INVXL U24392 ( .A(conv_3[282]), .Y(n32603) );
  INVXL U24393 ( .A(conv_3[327]), .Y(n33282) );
  OAI22XL U24394 ( .A0(n16668), .A1(n32603), .B0(n18321), .B1(n33282), .Y(
        n19554) );
  AOI211XL U24395 ( .A0(conv_3[297]), .A1(n22347), .B0(n19555), .C0(n19554), 
        .Y(n21434) );
  INVXL U24396 ( .A(conv_3[357]), .Y(n33728) );
  INVXL U24397 ( .A(conv_3[342]), .Y(n31986) );
  OAI22XL U24398 ( .A0(n19401), .A1(n33728), .B0(n22717), .B1(n31986), .Y(
        n19557) );
  INVXL U24399 ( .A(conv_3[372]), .Y(n31643) );
  INVXL U24400 ( .A(conv_3[387]), .Y(n34169) );
  OAI22XL U24401 ( .A0(n22612), .A1(n31643), .B0(n22716), .B1(n34169), .Y(
        n19556) );
  OAI22XL U24402 ( .A0(n21434), .A1(n26474), .B0(n21433), .B1(n26039), .Y(
        n19562) );
  INVXL U24403 ( .A(conv_3[207]), .Y(n31864) );
  INVXL U24404 ( .A(conv_3[177]), .Y(n31583) );
  INVXL U24405 ( .A(conv_3[162]), .Y(n32295) );
  OAI22XL U24406 ( .A0(n19902), .A1(n31583), .B0(n22717), .B1(n32295), .Y(
        n19559) );
  OAI22XL U24407 ( .A0(n25975), .A1(n21435), .B0(n21430), .B1(n35198), .Y(
        n19561) );
  AOI211XL U24408 ( .A0(n16755), .A1(n20568), .B0(n19562), .C0(n19561), .Y(
        n19563) );
  NAND4XL U24409 ( .A(n19566), .B(n19565), .C(n19564), .D(n19563), .Y(n19593)
         );
  INVXL U24410 ( .A(conv_3[238]), .Y(n33898) );
  AOI22XL U24411 ( .A0(n16666), .A1(conv_3[178]), .B0(n25299), .B1(conv_3[163]), .Y(n19567) );
  NAND2XL U24412 ( .A(n19568), .B(n19567), .Y(n21405) );
  AOI22XL U24413 ( .A0(n16660), .A1(n21405), .B0(n26081), .B1(n21410), .Y(
        n19589) );
  INVXL U24414 ( .A(conv_3[28]), .Y(n34414) );
  AOI22XL U24415 ( .A0(n21992), .A1(conv_3[13]), .B0(n21991), .B1(n21402), .Y(
        n19572) );
  INVXL U24416 ( .A(conv_3[448]), .Y(n32143) );
  OAI22XL U24417 ( .A0(n21810), .A1(n32143), .B0(n16669), .B1(n34003), .Y(
        n19569) );
  AOI211XL U24418 ( .A0(conv_3[433]), .A1(n22021), .B0(n19570), .C0(n19569), 
        .Y(n19571) );
  OAI211XL U24419 ( .A0(n34414), .A1(n21953), .B0(n19572), .C0(n19571), .Y(
        n20557) );
  INVXL U24420 ( .A(conv_3[58]), .Y(n34160) );
  INVXL U24421 ( .A(conv_3[43]), .Y(n31297) );
  INVXL U24422 ( .A(conv_3[88]), .Y(n32150) );
  OAI22XL U24423 ( .A0(n22717), .A1(n31297), .B0(n18321), .B1(n32150), .Y(
        n19573) );
  AOI22XL U24424 ( .A0(conv_3[223]), .A1(n26082), .B0(n26276), .B1(n21418), 
        .Y(n19577) );
  INVXL U24425 ( .A(N17708), .Y(n22713) );
  NAND2XL U24426 ( .A(n22713), .B(n21402), .Y(n20550) );
  INVXL U24427 ( .A(n20554), .Y(n21403) );
  OAI2BB1XL U24428 ( .A0N(n20550), .A1N(n19575), .B0(n28528), .Y(n19576) );
  OAI211XL U24429 ( .A0(n21408), .A1(n35239), .B0(n19577), .C0(n19576), .Y(
        n19587) );
  INVXL U24430 ( .A(conv_3[343]), .Y(n32213) );
  OAI22XL U24431 ( .A0(n22612), .A1(n32121), .B0(n22717), .B1(n32213), .Y(
        n19579) );
  INVXL U24432 ( .A(conv_3[358]), .Y(n34749) );
  OAI22XL U24433 ( .A0(n19902), .A1(n34749), .B0(n18750), .B1(n34142), .Y(
        n19578) );
  AOI22XL U24434 ( .A0(n16666), .A1(conv_3[118]), .B0(n16662), .B1(conv_3[133]), .Y(n19581) );
  NAND2XL U24435 ( .A(n19581), .B(n19580), .Y(n21404) );
  AOI22XL U24436 ( .A0(n35236), .A1(n21404), .B0(n35231), .B1(n21409), .Y(
        n19585) );
  AOI22XL U24437 ( .A0(n16716), .A1(conv_3[313]), .B0(n22690), .B1(conv_3[283]), .Y(n19582) );
  NAND2XL U24438 ( .A(n19583), .B(n19582), .Y(n21411) );
  NAND2XL U24439 ( .A(n16671), .B(n21411), .Y(n19584) );
  OAI211XL U24440 ( .A0(n21407), .A1(n26039), .B0(n19585), .C0(n19584), .Y(
        n19586) );
  AOI211XL U24441 ( .A0(n16755), .A1(n20557), .B0(n19587), .C0(n19586), .Y(
        n19588) );
  OAI211XL U24442 ( .A0(n33898), .A1(n26085), .B0(n19589), .C0(n19588), .Y(
        n19592) );
  NOR3XL U24443 ( .A(pool[129]), .B(n19593), .C(n19592), .Y(n19603) );
  NOR4BBXL U24444 ( .AN(n19593), .BN(n19592), .C(n19591), .D(n19590), .Y(
        n19599) );
  OR2XL U24445 ( .A(n19742), .B(n19741), .Y(n19594) );
  NOR4XL U24446 ( .A(n19597), .B(n19596), .C(n19595), .D(n19594), .Y(n19598)
         );
  NAND4BBXL U24447 ( .AN(n19601), .BN(n19600), .C(n19599), .D(n19598), .Y(
        n19602) );
  NAND2XL U24448 ( .A(n35026), .B(pool[125]), .Y(n19607) );
  OAI21XL U24449 ( .A0(n19608), .A1(n35026), .B0(n19607), .Y(N29341) );
  MXI2XL U24450 ( .A(n19626), .B(n19629), .S0(n19689), .Y(n19609) );
  OAI32XL U24451 ( .A0(n18010), .A1(n19694), .A2(n19629), .B0(n19609), .B1(
        n19630), .Y(n19618) );
  AOI221XL U24452 ( .A0(n19612), .A1(n19698), .B0(n19622), .B1(n19611), .C0(
        n19613), .Y(n19621) );
  AOI22XL U24453 ( .A0(n19614), .A1(n19652), .B0(n19698), .B1(n19613), .Y(
        n19615) );
  OAI22XL U24454 ( .A0(n19622), .A1(n19617), .B0(n19616), .B1(n19615), .Y(
        n19620) );
  ADDHXL U24455 ( .A(affine_2[19]), .B(n19618), .CO(DP_OP_5170J1_126_4278_n67), 
        .S(n19619) );
  ADDFX1 U24456 ( .A(n19621), .B(n19620), .CI(n19619), .CO(n20103), .S(n19681)
         );
  MXI2XL U24457 ( .A(n19626), .B(n19629), .S0(n19694), .Y(n19623) );
  OAI32XL U24458 ( .A0(n18010), .A1(n19666), .A2(n19629), .B0(n19623), .B1(
        n19630), .Y(n19624) );
  ADDFX1 U24459 ( .A(n19625), .B(affine_2[18]), .CI(n19624), .CO(n19680), .S(
        n19738) );
  NAND2XL U24460 ( .A(n19626), .B(n19630), .Y(n19628) );
  MXI2XL U24461 ( .A(n19626), .B(n19629), .S0(n19666), .Y(n19627) );
  OAI22XL U24462 ( .A0(n19698), .A1(n19628), .B0(n19627), .B1(n19630), .Y(
        n19631) );
  AOI21XL U24463 ( .A0(n19698), .A1(n18010), .B0(n19629), .Y(n19658) );
  ADDHXL U24464 ( .A(affine_2[17]), .B(n19631), .CO(n19737), .S(n19656) );
  AOI222XL U24465 ( .A0(n33367), .A1(affine_2[20]), .B0(n16674), .B1(n19633), 
        .C0(weight_2_bias_2[4]), .C1(n20614), .Y(n19634) );
  INVXL U24466 ( .A(n19634), .Y(n16541) );
  MXI2XL U24467 ( .A(n19647), .B(n19650), .S0(n19689), .Y(n19635) );
  OAI32XL U24468 ( .A0(n17929), .A1(n19694), .A2(n19650), .B0(n19635), .B1(
        n19651), .Y(n19642) );
  AOI221XL U24469 ( .A0(n19637), .A1(n19698), .B0(n19643), .B1(n19636), .C0(
        n19638), .Y(n19730) );
  AOI22XL U24470 ( .A0(n17962), .A1(n19652), .B0(n19698), .B1(n19638), .Y(
        n19639) );
  ADDHXL U24471 ( .A(affine_2[35]), .B(n19642), .CO(DP_OP_5169J1_125_4278_n67), 
        .S(n19728) );
  MXI2XL U24472 ( .A(n19647), .B(n19650), .S0(n19694), .Y(n19644) );
  OAI32XL U24473 ( .A0(n17929), .A1(n19666), .A2(n19650), .B0(n19644), .B1(
        n19651), .Y(n19645) );
  ADDFX1 U24474 ( .A(n19646), .B(affine_2[34]), .CI(n19645), .CO(n19732), .S(
        n19686) );
  NAND2XL U24475 ( .A(n19647), .B(n19651), .Y(n19649) );
  MXI2XL U24476 ( .A(n19647), .B(n19650), .S0(n19666), .Y(n19648) );
  OAI22XL U24477 ( .A0(n19698), .A1(n19649), .B0(n19648), .B1(n19651), .Y(
        n19653) );
  AOI21XL U24478 ( .A0(n19698), .A1(n17929), .B0(n19650), .Y(n19725) );
  NOR2XL U24479 ( .A(n19652), .B(n19651), .Y(n19720) );
  ADDHXL U24480 ( .A(affine_2[33]), .B(n19653), .CO(n19685), .S(n19723) );
  AOI222XL U24481 ( .A0(n33367), .A1(affine_2[35]), .B0(n16674), .B1(n19654), 
        .C0(weight_2_bias_3[3]), .C1(n20614), .Y(n19655) );
  INVXL U24482 ( .A(n19655), .Y(n16558) );
  ADDFX1 U24483 ( .A(n19658), .B(n19657), .CI(n19656), .CO(n19736), .S(n19659)
         );
  AOI222XL U24484 ( .A0(n33367), .A1(affine_2[17]), .B0(n16674), .B1(n19659), 
        .C0(weight_2_bias_2[1]), .C1(n20614), .Y(n19660) );
  INVXL U24485 ( .A(n19660), .Y(n16544) );
  AOI21XL U24486 ( .A0(n19698), .A1(n18078), .B0(n19693), .Y(n19670) );
  NAND2XL U24487 ( .A(n18084), .B(n19691), .Y(n19662) );
  MXI2XL U24488 ( .A(n18084), .B(n19693), .S0(n19666), .Y(n19661) );
  OAI22XL U24489 ( .A0(n19698), .A1(n19662), .B0(n19661), .B1(n19691), .Y(
        n19667) );
  AOI222XL U24490 ( .A0(n33367), .A1(affine_2[1]), .B0(n16674), .B1(n19663), 
        .C0(weight_2_bias_1[1]), .C1(n20614), .Y(n19664) );
  INVXL U24491 ( .A(n19664), .Y(n16578) );
  MXI2XL U24492 ( .A(n18084), .B(n19693), .S0(n19694), .Y(n19665) );
  OAI32XL U24493 ( .A0(n18078), .A1(n19666), .A2(n19693), .B0(n19665), .B1(
        n19691), .Y(n19708) );
  ADDHXL U24494 ( .A(affine_2[1]), .B(n19667), .CO(n19711), .S(n19668) );
  ADDFX1 U24495 ( .A(n19670), .B(n19669), .CI(n19668), .CO(n19710), .S(n19663)
         );
  AOI222XL U24496 ( .A0(n33367), .A1(affine_2[2]), .B0(n16674), .B1(n19671), 
        .C0(weight_2_bias_1[2]), .C1(n20614), .Y(n19672) );
  INVXL U24497 ( .A(n19672), .Y(n16577) );
  ADDHXL U24498 ( .A(affine_2[16]), .B(n19673), .CO(n19657), .S(n19674) );
  AOI222XL U24499 ( .A0(n33367), .A1(affine_2[16]), .B0(n16674), .B1(n19674), 
        .C0(weight_2_bias_2[0]), .C1(n20614), .Y(n19675) );
  INVXL U24500 ( .A(n19675), .Y(n16545) );
  ADDHXL U24501 ( .A(affine_2[0]), .B(n19676), .CO(n19669), .S(n19677) );
  AOI222XL U24502 ( .A0(n33367), .A1(affine_2[0]), .B0(n16674), .B1(n19677), 
        .C0(weight_2_bias_1[0]), .C1(n20614), .Y(n19678) );
  INVXL U24503 ( .A(n19678), .Y(n16579) );
  ADDFX1 U24504 ( .A(n19681), .B(n19680), .CI(n19679), .CO(n20102), .S(n19682)
         );
  AOI222XL U24505 ( .A0(n33367), .A1(affine_2[19]), .B0(n16674), .B1(n19682), 
        .C0(weight_2_bias_2[3]), .C1(n20614), .Y(n19683) );
  INVXL U24506 ( .A(n19683), .Y(n16542) );
  ADDFX1 U24507 ( .A(n19686), .B(n19685), .CI(n19684), .CO(n19731), .S(n19687)
         );
  AOI222XL U24508 ( .A0(n33367), .A1(affine_2[34]), .B0(n16674), .B1(n19687), 
        .C0(weight_2_bias_3[2]), .C1(n20614), .Y(n19688) );
  INVXL U24509 ( .A(n19688), .Y(n16559) );
  MXI2XL U24510 ( .A(n18084), .B(n19693), .S0(n19689), .Y(n19692) );
  OAI32XL U24511 ( .A0(n18078), .A1(n19694), .A2(n19693), .B0(n19692), .B1(
        n19691), .Y(n19704) );
  AOI221XL U24512 ( .A0(n19696), .A1(n19698), .B0(n19703), .B1(n19695), .C0(
        n19697), .Y(n19707) );
  AOI22XL U24513 ( .A0(n18106), .A1(n19652), .B0(n19698), .B1(n19697), .Y(
        n19700) );
  OAI22XL U24514 ( .A0(n19703), .A1(n19702), .B0(n19701), .B1(n19700), .Y(
        n19706) );
  ADDHXL U24515 ( .A(affine_2[3]), .B(n19704), .CO(DP_OP_5171J1_127_4278_n67), 
        .S(n19705) );
  ADDFX1 U24516 ( .A(n19707), .B(n19706), .CI(n19705), .CO(n20116), .S(n19717)
         );
  ADDFX1 U24517 ( .A(n19712), .B(n19711), .CI(n19710), .CO(n19715), .S(n19671)
         );
  AOI222XL U24518 ( .A0(n33367), .A1(affine_2[4]), .B0(n16674), .B1(n19713), 
        .C0(weight_2_bias_1[4]), .C1(n20614), .Y(n19714) );
  INVXL U24519 ( .A(n19714), .Y(n16575) );
  ADDFX1 U24520 ( .A(n19717), .B(n19716), .CI(n19715), .CO(n20115), .S(n19718)
         );
  AOI222XL U24521 ( .A0(n33367), .A1(affine_2[3]), .B0(n16674), .B1(n19718), 
        .C0(weight_2_bias_1[3]), .C1(n20614), .Y(n19719) );
  INVXL U24522 ( .A(n19719), .Y(n16576) );
  ADDHXL U24523 ( .A(affine_2[32]), .B(n19720), .CO(n19724), .S(n19721) );
  AOI222XL U24524 ( .A0(n33367), .A1(affine_2[32]), .B0(n16674), .B1(n19721), 
        .C0(weight_2_bias_3[0]), .C1(n20614), .Y(n19722) );
  INVXL U24525 ( .A(n19722), .Y(n16561) );
  ADDFX1 U24526 ( .A(n19725), .B(n19724), .CI(n19723), .CO(n19684), .S(n19726)
         );
  AOI222XL U24527 ( .A0(n33367), .A1(affine_2[33]), .B0(n16674), .B1(n19726), 
        .C0(weight_2_bias_3[1]), .C1(n20614), .Y(n19727) );
  INVXL U24528 ( .A(n19727), .Y(n16560) );
  ADDFX1 U24529 ( .A(n19730), .B(n19729), .CI(n19728), .CO(n20123), .S(n19733)
         );
  ADDFX1 U24530 ( .A(n19733), .B(n19732), .CI(n19731), .CO(n20122), .S(n19654)
         );
  AOI222XL U24531 ( .A0(n33367), .A1(affine_2[36]), .B0(n16674), .B1(n19734), 
        .C0(weight_2_bias_3[4]), .C1(n20614), .Y(n19735) );
  INVXL U24532 ( .A(n19735), .Y(n16557) );
  ADDFX1 U24533 ( .A(n19738), .B(n19737), .CI(n19736), .CO(n19679), .S(n19739)
         );
  AOI222XL U24534 ( .A0(n33367), .A1(affine_2[18]), .B0(n16674), .B1(n19739), 
        .C0(weight_2_bias_2[2]), .C1(n20614), .Y(n19740) );
  INVXL U24535 ( .A(n19740), .Y(n16543) );
  AOI22XL U24536 ( .A0(n35026), .A1(n19742), .B0(n19741), .B1(n35027), .Y(
        N29345) );
  AOI22XL U24537 ( .A0(n16734), .A1(conv_1[405]), .B0(n21954), .B1(conv_1[390]), .Y(n19746) );
  INVXL U24538 ( .A(conv_1[465]), .Y(n33510) );
  INVXL U24539 ( .A(conv_1[450]), .Y(n27424) );
  AOI22XL U24540 ( .A0(n20735), .A1(n33510), .B0(n27424), .B1(n18634), .Y(
        n25297) );
  AOI22XL U24541 ( .A0(n21990), .A1(conv_1[420]), .B0(n21991), .B1(n25297), 
        .Y(n19745) );
  AOI22XL U24542 ( .A0(conv_1[15]), .A1(n22015), .B0(n21887), .B1(conv_1[435]), 
        .Y(n19744) );
  NAND2XL U24543 ( .A(conv_1[0]), .B(n21992), .Y(n19743) );
  NAND4XL U24544 ( .A(n19746), .B(n19745), .C(n19744), .D(n19743), .Y(n20193)
         );
  INVXL U24545 ( .A(conv_1[255]), .Y(n33526) );
  INVXL U24546 ( .A(conv_1[240]), .Y(n33536) );
  AOI22XL U24547 ( .A0(n20735), .A1(n33526), .B0(n33536), .B1(n18634), .Y(
        n25298) );
  INVXL U24548 ( .A(conv_1[225]), .Y(n33875) );
  INVXL U24549 ( .A(conv_1[210]), .Y(n33871) );
  AOI22XL U24550 ( .A0(n20735), .A1(n33875), .B0(n33871), .B1(n18634), .Y(
        n25294) );
  INVXL U24551 ( .A(N17708), .Y(n22743) );
  AOI22XL U24552 ( .A0(n20735), .A1(conv_1[495]), .B0(conv_1[480]), .B1(n19253), .Y(n25304) );
  INVXL U24553 ( .A(n25304), .Y(n21465) );
  AOI22XL U24554 ( .A0(n34952), .A1(n25297), .B0(n34950), .B1(n21465), .Y(
        n19750) );
  AOI22XL U24555 ( .A0(n22762), .A1(conv_1[165]), .B0(n16662), .B1(conv_1[180]), .Y(n19748) );
  AOI22XL U24556 ( .A0(n22759), .A1(conv_1[150]), .B0(n16673), .B1(conv_1[195]), .Y(n19747) );
  NAND2XL U24557 ( .A(n19748), .B(n19747), .Y(n21460) );
  AOI22XL U24558 ( .A0(n20735), .A1(conv_1[525]), .B0(conv_1[510]), .B1(n19253), .Y(n25305) );
  AOI22XL U24559 ( .A0(n16667), .A1(n21460), .B0(n34954), .B1(n21468), .Y(
        n19749) );
  OAI211XL U24560 ( .A0(n21466), .A1(n34958), .B0(n19750), .C0(n19749), .Y(
        n19762) );
  AOI22XL U24561 ( .A0(n21831), .A1(n25298), .B0(n21468), .B1(n21830), .Y(
        n20190) );
  AOI22XL U24562 ( .A0(n25299), .A1(conv_1[30]), .B0(n16673), .B1(conv_1[75]), 
        .Y(n19752) );
  AOI22XL U24563 ( .A0(n22762), .A1(conv_1[45]), .B0(n16662), .B1(conv_1[60]), 
        .Y(n19751) );
  NAND2XL U24564 ( .A(n19752), .B(n19751), .Y(n21467) );
  AOI22XL U24565 ( .A0(n22762), .A1(conv_1[345]), .B0(n16673), .B1(conv_1[375]), .Y(n19754) );
  AOI22XL U24566 ( .A0(n16716), .A1(conv_1[360]), .B0(n22690), .B1(conv_1[330]), .Y(n19753) );
  AOI22XL U24567 ( .A0(n25299), .A1(conv_1[90]), .B0(n16673), .B1(conv_1[135]), 
        .Y(n19756) );
  AOI22XL U24568 ( .A0(n22762), .A1(conv_1[105]), .B0(n16662), .B1(conv_1[120]), .Y(n19755) );
  NAND2XL U24569 ( .A(n19756), .B(n19755), .Y(n21469) );
  INVX2 U24570 ( .A(n18196), .Y(n34961) );
  AOI22XL U24571 ( .A0(n16716), .A1(conv_1[300]), .B0(n18658), .B1(conv_1[270]), .Y(n19758) );
  AOI22XL U24572 ( .A0(n22762), .A1(conv_1[285]), .B0(n16673), .B1(conv_1[315]), .Y(n19757) );
  NAND2XL U24573 ( .A(n19758), .B(n19757), .Y(n21459) );
  AOI22XL U24574 ( .A0(n28528), .A1(n21469), .B0(n34961), .B1(n21459), .Y(
        n19759) );
  OAI211XL U24575 ( .A0(n20190), .A1(n34969), .B0(n19760), .C0(n19759), .Y(
        n19761) );
  AOI211XL U24576 ( .A0(n28465), .A1(n20193), .B0(n19762), .C0(n19761), .Y(
        n20101) );
  INVXL U24577 ( .A(conv_1[464]), .Y(n28754) );
  AOI22XL U24578 ( .A0(n20735), .A1(n28738), .B0(n28754), .B1(n18516), .Y(
        n22722) );
  AOI22XL U24579 ( .A0(conv_1[239]), .A1(n21999), .B0(n34952), .B1(n22722), 
        .Y(n19785) );
  AOI22XL U24580 ( .A0(n22762), .A1(conv_1[119]), .B0(n16673), .B1(conv_1[149]), .Y(n19764) );
  AOI22XL U24581 ( .A0(n18810), .A1(conv_1[134]), .B0(n22759), .B1(conv_1[104]), .Y(n19763) );
  NAND2XL U24582 ( .A(n19764), .B(n19763), .Y(n21709) );
  AOI22XL U24583 ( .A0(n22616), .A1(conv_1[284]), .B0(n16673), .B1(conv_1[329]), .Y(n19766) );
  AOI22XL U24584 ( .A0(n22762), .A1(conv_1[299]), .B0(n16662), .B1(conv_1[314]), .Y(n19765) );
  NAND2XL U24585 ( .A(n19766), .B(n19765), .Y(n21707) );
  AOI22XL U24586 ( .A0(n28528), .A1(n21709), .B0(n34961), .B1(n21707), .Y(
        n19784) );
  AOI22XL U24587 ( .A0(n20735), .A1(conv_1[509]), .B0(conv_1[494]), .B1(n18526), .Y(n22720) );
  AOI22XL U24588 ( .A0(n20735), .A1(conv_1[539]), .B0(conv_1[524]), .B1(n18516), .Y(n22721) );
  INVXL U24589 ( .A(conv_1[59]), .Y(n33054) );
  INVXL U24590 ( .A(conv_1[74]), .Y(n27211) );
  INVXL U24591 ( .A(conv_1[89]), .Y(n26838) );
  OAI22XL U24592 ( .A0(n22612), .A1(n27211), .B0(n24039), .B1(n26838), .Y(
        n19768) );
  AOI211XL U24593 ( .A0(conv_1[44]), .A1(n22616), .B0(n19769), .C0(n19768), 
        .Y(n21724) );
  INVXL U24594 ( .A(conv_1[194]), .Y(n32995) );
  INVXL U24595 ( .A(conv_1[164]), .Y(n23375) );
  INVXL U24596 ( .A(conv_1[209]), .Y(n33122) );
  OAI22XL U24597 ( .A0(n16668), .A1(n23375), .B0(n22716), .B1(n33122), .Y(
        n19770) );
  INVXL U24598 ( .A(conv_1[374]), .Y(n33134) );
  INVXL U24599 ( .A(conv_1[359]), .Y(n28820) );
  INVXL U24600 ( .A(conv_1[344]), .Y(n28828) );
  OAI22XL U24601 ( .A0(n19902), .A1(n28820), .B0(n22717), .B1(n28828), .Y(
        n19772) );
  AOI211XL U24602 ( .A0(conv_1[389]), .A1(n16673), .B0(n19773), .C0(n19772), 
        .Y(n21705) );
  OAI22XL U24603 ( .A0(n21713), .A1(n28577), .B0(n21705), .B1(n35196), .Y(
        n19774) );
  AOI211XL U24604 ( .A0(n21708), .A1(n24056), .B0(n19775), .C0(n19774), .Y(
        n19783) );
  AOI22XL U24605 ( .A0(n21990), .A1(conv_1[434]), .B0(n16734), .B1(conv_1[419]), .Y(n19779) );
  AOI22XL U24606 ( .A0(n21954), .A1(conv_1[404]), .B0(n21991), .B1(n22722), 
        .Y(n19778) );
  AOI22XL U24607 ( .A0(conv_1[29]), .A1(n22015), .B0(n21887), .B1(conv_1[449]), 
        .Y(n19777) );
  NAND2XL U24608 ( .A(conv_1[14]), .B(n21992), .Y(n19776) );
  NAND4XL U24609 ( .A(n19779), .B(n19778), .C(n19777), .D(n19776), .Y(n20201)
         );
  INVXL U24610 ( .A(conv_1[224]), .Y(n28606) );
  OAI22XL U24611 ( .A0(n22721), .A1(n21959), .B0(n28606), .B1(n22030), .Y(
        n19781) );
  AOI22XL U24612 ( .A0(n20735), .A1(conv_1[269]), .B0(conv_1[254]), .B1(n18634), .Y(n22712) );
  OAI22XL U24613 ( .A0(n22720), .A1(n21960), .B0(n22712), .B1(n20491), .Y(
        n19780) );
  AOI211XL U24614 ( .A0(n28465), .A1(n20201), .B0(n19781), .C0(n19780), .Y(
        n19782) );
  NAND4XL U24615 ( .A(n19785), .B(n19784), .C(n19783), .D(n19782), .Y(n20098)
         );
  INVXL U24616 ( .A(conv_1[468]), .Y(n26956) );
  INVXL U24617 ( .A(conv_1[453]), .Y(n27254) );
  AOI22XL U24618 ( .A0(n20735), .A1(n26956), .B0(n27254), .B1(n18634), .Y(
        n22635) );
  AOI22XL U24619 ( .A0(n21954), .A1(conv_1[393]), .B0(n21991), .B1(n22635), 
        .Y(n19789) );
  AOI22XL U24620 ( .A0(n21990), .A1(conv_1[423]), .B0(n21887), .B1(conv_1[438]), .Y(n19788) );
  AOI22XL U24621 ( .A0(conv_1[18]), .A1(n22015), .B0(n16734), .B1(conv_1[408]), 
        .Y(n19787) );
  NAND2XL U24622 ( .A(conv_1[3]), .B(n21992), .Y(n19786) );
  NAND4XL U24623 ( .A(n19789), .B(n19788), .C(n19787), .D(n19786), .Y(n20214)
         );
  INVXL U24624 ( .A(conv_1[228]), .Y(n23368) );
  INVXL U24625 ( .A(conv_1[528]), .Y(n32869) );
  INVXL U24626 ( .A(conv_1[513]), .Y(n30459) );
  AOI22XL U24627 ( .A0(n20735), .A1(n32869), .B0(n30459), .B1(n18634), .Y(
        n22644) );
  INVXL U24628 ( .A(conv_1[258]), .Y(n23472) );
  AOI22XL U24629 ( .A0(n21998), .A1(n22644), .B0(n22011), .B1(n22638), .Y(
        n19791) );
  INVXL U24630 ( .A(conv_1[498]), .Y(n29546) );
  INVXL U24631 ( .A(conv_1[483]), .Y(n27229) );
  AOI22XL U24632 ( .A0(n20735), .A1(n29546), .B0(n27229), .B1(n18516), .Y(
        n22643) );
  NAND2XL U24633 ( .A(n34950), .B(n22643), .Y(n19790) );
  OAI211XL U24634 ( .A0(n22008), .A1(n23368), .B0(n19791), .C0(n19790), .Y(
        n19807) );
  AOI22XL U24635 ( .A0(n16744), .A1(conv_1[213]), .B0(n34952), .B1(n22635), 
        .Y(n19805) );
  INVX2 U24636 ( .A(n28479), .Y(n28528) );
  AOI22XL U24637 ( .A0(n25299), .A1(conv_1[93]), .B0(n16673), .B1(conv_1[138]), 
        .Y(n19793) );
  AOI22XL U24638 ( .A0(n22762), .A1(conv_1[108]), .B0(n16662), .B1(conv_1[123]), .Y(n19792) );
  NAND2XL U24639 ( .A(n19793), .B(n19792), .Y(n21482) );
  AOI22XL U24640 ( .A0(n16716), .A1(conv_1[183]), .B0(n16673), .B1(conv_1[198]), .Y(n19795) );
  AOI22XL U24641 ( .A0(n22762), .A1(conv_1[168]), .B0(n22759), .B1(conv_1[153]), .Y(n19794) );
  NAND2XL U24642 ( .A(n19795), .B(n19794), .Y(n21483) );
  AOI22XL U24643 ( .A0(n28528), .A1(n21482), .B0(n16667), .B1(n21483), .Y(
        n19804) );
  AOI22XL U24644 ( .A0(n22616), .A1(conv_1[333]), .B0(n16673), .B1(conv_1[378]), .Y(n19797) );
  NAND2XL U24645 ( .A(n19797), .B(n19796), .Y(n21481) );
  NAND2XL U24646 ( .A(n21688), .B(n22644), .Y(n20207) );
  NAND2XL U24647 ( .A(n20206), .B(n20207), .Y(n21485) );
  AOI22XL U24648 ( .A0(n35234), .A1(n21481), .B0(n21485), .B1(n24056), .Y(
        n19803) );
  AOI22XL U24649 ( .A0(n20978), .A1(conv_1[48]), .B0(n16673), .B1(conv_1[78]), 
        .Y(n19799) );
  AOI22XL U24650 ( .A0(n16716), .A1(conv_1[63]), .B0(n22690), .B1(conv_1[33]), 
        .Y(n19798) );
  NAND2XL U24651 ( .A(n19799), .B(n19798), .Y(n21480) );
  AOI22XL U24652 ( .A0(n22690), .A1(conv_1[273]), .B0(n16673), .B1(conv_1[318]), .Y(n19801) );
  NAND2XL U24653 ( .A(n19801), .B(n19800), .Y(n21484) );
  NAND4XL U24654 ( .A(n19805), .B(n19804), .C(n19803), .D(n19802), .Y(n19806)
         );
  INVXL U24655 ( .A(conv_1[467]), .Y(n26989) );
  INVXL U24656 ( .A(conv_1[452]), .Y(n27384) );
  AOI22XL U24657 ( .A0(n20735), .A1(n26989), .B0(n27384), .B1(n19253), .Y(
        n22662) );
  AOI22XL U24658 ( .A0(n16734), .A1(conv_1[407]), .B0(n21991), .B1(n22662), 
        .Y(n19811) );
  AOI22XL U24659 ( .A0(n21990), .A1(conv_1[422]), .B0(n21954), .B1(conv_1[392]), .Y(n19810) );
  AOI22XL U24660 ( .A0(n21887), .A1(conv_1[437]), .B0(conv_1[2]), .B1(n21992), 
        .Y(n19809) );
  NAND2XL U24661 ( .A(conv_1[17]), .B(n22015), .Y(n19808) );
  NAND4XL U24662 ( .A(n19811), .B(n19810), .C(n19809), .D(n19808), .Y(n20230)
         );
  INVXL U24663 ( .A(conv_1[527]), .Y(n30465) );
  INVXL U24664 ( .A(conv_1[512]), .Y(n26985) );
  AOI22XL U24665 ( .A0(n20735), .A1(n30465), .B0(n26985), .B1(n19253), .Y(
        n22657) );
  INVXL U24666 ( .A(conv_1[497]), .Y(n23421) );
  INVXL U24667 ( .A(conv_1[482]), .Y(n27378) );
  AOI22XL U24668 ( .A0(n20735), .A1(n23421), .B0(n27378), .B1(n18634), .Y(
        n22656) );
  AND2XL U24669 ( .A(n36246), .B(n22656), .Y(n21517) );
  AOI21XL U24670 ( .A0(n22765), .A1(n22657), .B0(n21517), .Y(n20227) );
  INVXL U24671 ( .A(n20227), .Y(n21520) );
  NAND2XL U24672 ( .A(n21830), .B(n21520), .Y(n20223) );
  INVXL U24673 ( .A(N17708), .Y(n22765) );
  INVXL U24674 ( .A(conv_1[257]), .Y(n23968) );
  INVXL U24675 ( .A(conv_1[242]), .Y(n24387) );
  AOI22XL U24676 ( .A0(n20735), .A1(n23968), .B0(n24387), .B1(n18526), .Y(
        n22655) );
  AOI22XL U24677 ( .A0(n34952), .A1(n22662), .B0(n21833), .B1(n22655), .Y(
        n19812) );
  NAND2XL U24678 ( .A(n21831), .B(n22655), .Y(n20224) );
  AOI32XL U24679 ( .A0(n20223), .A1(n19812), .A2(n20224), .B0(n34969), .B1(
        n19812), .Y(n19828) );
  AOI22XL U24680 ( .A0(n16744), .A1(conv_1[212]), .B0(n34950), .B1(n22656), 
        .Y(n19826) );
  AOI22XL U24681 ( .A0(n16716), .A1(conv_1[362]), .B0(n16673), .B1(conv_1[377]), .Y(n19813) );
  NAND2XL U24682 ( .A(n19814), .B(n19813), .Y(n21515) );
  AOI22XL U24683 ( .A0(conv_1[227]), .A1(n21999), .B0(n35234), .B1(n21515), 
        .Y(n19825) );
  AOI22XL U24684 ( .A0(n16716), .A1(conv_1[62]), .B0(n16673), .B1(conv_1[77]), 
        .Y(n19816) );
  NAND2XL U24685 ( .A(n19816), .B(n19815), .Y(n21516) );
  AOI22XL U24686 ( .A0(n25299), .A1(conv_1[272]), .B0(n16673), .B1(conv_1[317]), .Y(n19817) );
  NAND2XL U24687 ( .A(n19818), .B(n19817), .Y(n21521) );
  AOI22XL U24688 ( .A0(n16716), .A1(conv_1[122]), .B0(n16673), .B1(conv_1[137]), .Y(n19820) );
  NAND2XL U24689 ( .A(n19820), .B(n19819), .Y(n21519) );
  AOI22XL U24690 ( .A0(n22690), .A1(conv_1[152]), .B0(n16673), .B1(conv_1[197]), .Y(n19821) );
  NAND2XL U24691 ( .A(n19822), .B(n19821), .Y(n21522) );
  AOI22XL U24692 ( .A0(n28528), .A1(n21519), .B0(n16667), .B1(n21522), .Y(
        n19823) );
  NAND4XL U24693 ( .A(n19826), .B(n19825), .C(n19824), .D(n19823), .Y(n19827)
         );
  INVXL U24694 ( .A(conv_1[466]), .Y(n27015) );
  INVXL U24695 ( .A(conv_1[451]), .Y(n27437) );
  AOI22XL U24696 ( .A0(n35269), .A1(n27015), .B0(n27437), .B1(n18634), .Y(
        n22693) );
  AOI22XL U24697 ( .A0(n16734), .A1(conv_1[406]), .B0(n21991), .B1(n22693), 
        .Y(n19833) );
  AOI22XL U24698 ( .A0(n21990), .A1(conv_1[421]), .B0(n21887), .B1(conv_1[436]), .Y(n19832) );
  AOI22XL U24699 ( .A0(conv_1[16]), .A1(n22015), .B0(n21954), .B1(conv_1[391]), 
        .Y(n19831) );
  NAND2XL U24700 ( .A(conv_1[1]), .B(n21992), .Y(n19830) );
  NAND4XL U24701 ( .A(n19833), .B(n19832), .C(n19831), .D(n19830), .Y(n20218)
         );
  AOI22XL U24702 ( .A0(n20735), .A1(conv_1[496]), .B0(conv_1[481]), .B1(n18526), .Y(n22682) );
  AOI22XL U24703 ( .A0(n20735), .A1(conv_1[526]), .B0(conv_1[511]), .B1(n18526), .Y(n22683) );
  AOI22XL U24704 ( .A0(n35236), .A1(n19834), .B0(conv_1[211]), .B1(n16744), 
        .Y(n19836) );
  INVXL U24705 ( .A(conv_1[256]), .Y(n21798) );
  INVXL U24706 ( .A(conv_1[241]), .Y(n24437) );
  AOI22XL U24707 ( .A0(n20735), .A1(n21798), .B0(n24437), .B1(n18526), .Y(
        n22696) );
  NAND2XL U24708 ( .A(n22011), .B(n22696), .Y(n19835) );
  OAI211XL U24709 ( .A0(n22682), .A1(n21960), .B0(n19836), .C0(n19835), .Y(
        n19852) );
  AOI22XL U24710 ( .A0(n16716), .A1(conv_1[121]), .B0(n18658), .B1(conv_1[91]), 
        .Y(n19837) );
  AND2XL U24711 ( .A(n19838), .B(n19837), .Y(n21503) );
  NAND2XL U24712 ( .A(n22713), .B(n22693), .Y(n21496) );
  OAI22XL U24713 ( .A0(n21503), .A1(n28479), .B0(n26274), .B1(n21496), .Y(
        n19850) );
  INVXL U24714 ( .A(conv_1[76]), .Y(n27029) );
  INVXL U24715 ( .A(conv_1[46]), .Y(n27471) );
  INVXL U24716 ( .A(conv_1[31]), .Y(n24678) );
  OAI22XL U24717 ( .A0(n22546), .A1(n27471), .B0(n22550), .B1(n24678), .Y(
        n19839) );
  AOI22XL U24718 ( .A0(n16716), .A1(conv_1[181]), .B0(n22690), .B1(conv_1[151]), .Y(n19842) );
  AND2XL U24719 ( .A(n19842), .B(n19841), .Y(n21504) );
  OAI22XL U24720 ( .A0(n21497), .A1(n28575), .B0(n21504), .B1(n28577), .Y(
        n19849) );
  AOI22XL U24721 ( .A0(n22690), .A1(conv_1[271]), .B0(n16673), .B1(conv_1[316]), .Y(n19843) );
  NAND2XL U24722 ( .A(n19844), .B(n19843), .Y(n21506) );
  AOI22XL U24723 ( .A0(n34961), .A1(n21506), .B0(conv_1[226]), .B1(n21999), 
        .Y(n19848) );
  AOI22XL U24724 ( .A0(n35234), .A1(n21505), .B0(n21501), .B1(n24056), .Y(
        n19847) );
  NAND4BBXL U24725 ( .AN(n19850), .BN(n19849), .C(n19848), .D(n19847), .Y(
        n19851) );
  AOI222XL U24726 ( .A0(pool[5]), .A1(pool[6]), .B0(pool[5]), .B1(n34797), 
        .C0(pool[6]), .C1(n34797), .Y(n19853) );
  AOI222XL U24727 ( .A0(n34801), .A1(n34799), .B0(n34801), .B1(n19853), .C0(
        n34799), .C1(n19853), .Y(n19854) );
  AOI222XL U24728 ( .A0(n20160), .A1(pool[8]), .B0(n20160), .B1(n19854), .C0(
        pool[8]), .C1(n19854), .Y(n20039) );
  INVXL U24729 ( .A(conv_1[461]), .Y(n30029) );
  INVXL U24730 ( .A(conv_1[26]), .Y(n33201) );
  INVXL U24731 ( .A(conv_1[11]), .Y(n34553) );
  AOI22XL U24732 ( .A0(n21990), .A1(conv_1[431]), .B0(n16734), .B1(conv_1[416]), .Y(n19857) );
  AOI22XL U24733 ( .A0(n21887), .A1(conv_1[446]), .B0(n21954), .B1(conv_1[401]), .Y(n19856) );
  OAI211XL U24734 ( .A0(n34553), .A1(n22018), .B0(n19857), .C0(n19856), .Y(
        n19858) );
  AOI211XL U24735 ( .A0(n21991), .A1(n22590), .B0(n19859), .C0(n19858), .Y(
        n20287) );
  INVXL U24736 ( .A(conv_1[473]), .Y(n27177) );
  INVXL U24737 ( .A(conv_1[458]), .Y(n30041) );
  AOI22XL U24738 ( .A0(n20735), .A1(n27177), .B0(n30041), .B1(n19253), .Y(
        n22560) );
  AOI22XL U24739 ( .A0(n16734), .A1(conv_1[413]), .B0(n21991), .B1(n22560), 
        .Y(n19863) );
  AOI22XL U24740 ( .A0(n21887), .A1(conv_1[443]), .B0(n21954), .B1(conv_1[398]), .Y(n19862) );
  AOI22XL U24741 ( .A0(conv_1[23]), .A1(n22015), .B0(n21990), .B1(conv_1[428]), 
        .Y(n19861) );
  NAND2XL U24742 ( .A(conv_1[8]), .B(n21992), .Y(n19860) );
  NAND4XL U24743 ( .A(n19863), .B(n19862), .C(n19861), .D(n19860), .Y(n20281)
         );
  INVXL U24744 ( .A(conv_1[475]), .Y(n32890) );
  INVXL U24745 ( .A(conv_1[460]), .Y(n30048) );
  AOI22XL U24746 ( .A0(n20735), .A1(n32890), .B0(n30048), .B1(n18634), .Y(
        n22490) );
  AOI22XL U24747 ( .A0(n16734), .A1(conv_1[415]), .B0(n21991), .B1(n22490), 
        .Y(n19867) );
  AOI22XL U24748 ( .A0(n21887), .A1(conv_1[445]), .B0(n21954), .B1(conv_1[400]), .Y(n19866) );
  AOI22XL U24749 ( .A0(conv_1[25]), .A1(n22015), .B0(n21990), .B1(conv_1[430]), 
        .Y(n19865) );
  NAND2XL U24750 ( .A(conv_1[10]), .B(n21992), .Y(n19864) );
  NAND4XL U24751 ( .A(n19867), .B(n19866), .C(n19865), .D(n19864), .Y(n20297)
         );
  INVXL U24752 ( .A(conv_1[459]), .Y(n30035) );
  AOI22XL U24753 ( .A0(n20735), .A1(n26346), .B0(n30035), .B1(n18516), .Y(
        n22532) );
  AOI22XL U24754 ( .A0(n21954), .A1(conv_1[399]), .B0(n21991), .B1(n22532), 
        .Y(n19871) );
  AOI22XL U24755 ( .A0(n21990), .A1(conv_1[429]), .B0(n16734), .B1(conv_1[414]), .Y(n19870) );
  AOI22XL U24756 ( .A0(n21887), .A1(conv_1[444]), .B0(conv_1[9]), .B1(n21992), 
        .Y(n19869) );
  NAND2XL U24757 ( .A(conv_1[24]), .B(n22015), .Y(n19868) );
  NAND4XL U24758 ( .A(n19871), .B(n19870), .C(n19869), .D(n19868), .Y(n20306)
         );
  NOR4BXL U24759 ( .AN(n20287), .B(n20281), .C(n20297), .D(n20306), .Y(n20033)
         );
  AOI22XL U24760 ( .A0(n21990), .A1(conv_1[424]), .B0(n21887), .B1(conv_1[439]), .Y(n19875) );
  INVXL U24761 ( .A(conv_1[394]), .Y(n30764) );
  INVXL U24762 ( .A(conv_1[469]), .Y(n27011) );
  INVXL U24763 ( .A(conv_1[454]), .Y(n27397) );
  OAI22XL U24764 ( .A0(n18634), .A1(n27011), .B0(n27397), .B1(n35269), .Y(
        n22499) );
  OAI2BB2XL U24765 ( .B0(n16669), .B1(n30764), .A0N(n22499), .A1N(n21991), .Y(
        n19873) );
  INVXL U24766 ( .A(conv_1[19]), .Y(n27455) );
  INVXL U24767 ( .A(conv_1[409]), .Y(n35486) );
  OAI22XL U24768 ( .A0(n27455), .A1(n21953), .B0(n21944), .B1(n35486), .Y(
        n19872) );
  AOI211XL U24769 ( .A0(conv_1[4]), .A1(n21992), .B0(n19873), .C0(n19872), .Y(
        n19874) );
  NAND2XL U24770 ( .A(n19875), .B(n19874), .Y(n20245) );
  AOI22XL U24771 ( .A0(n20735), .A1(conv_1[259]), .B0(conv_1[244]), .B1(n18634), .Y(n22498) );
  INVXL U24772 ( .A(conv_1[514]), .Y(n27391) );
  AOI2BB2XL U24773 ( .B0(n27391), .B1(n19253), .A0N(n18634), .A1N(conv_1[529]), 
        .Y(n22510) );
  AOI22XL U24774 ( .A0(n34952), .A1(n22499), .B0(n21998), .B1(n22510), .Y(
        n19877) );
  NAND2XL U24775 ( .A(conv_1[229]), .B(n21999), .Y(n19876) );
  OAI211XL U24776 ( .A0(n22498), .A1(n20491), .B0(n19877), .C0(n19876), .Y(
        n19893) );
  INVXL U24777 ( .A(conv_1[499]), .Y(n30700) );
  INVXL U24778 ( .A(conv_1[484]), .Y(n27403) );
  AOI22XL U24779 ( .A0(n20735), .A1(n30700), .B0(n27403), .B1(n18634), .Y(
        n22509) );
  AOI22XL U24780 ( .A0(conv_1[214]), .A1(n16744), .B0(n34950), .B1(n22509), 
        .Y(n19891) );
  AOI22XL U24781 ( .A0(n20978), .A1(conv_1[49]), .B0(n16673), .B1(conv_1[79]), 
        .Y(n19879) );
  NAND2XL U24782 ( .A(n19879), .B(n19878), .Y(n21543) );
  NAND2XL U24783 ( .A(n22713), .B(n22510), .Y(n21538) );
  NAND2XL U24784 ( .A(n21535), .B(n21538), .Y(n21544) );
  AOI22XL U24785 ( .A0(n20978), .A1(conv_1[109]), .B0(n16673), .B1(conv_1[139]), .Y(n19880) );
  NAND2XL U24786 ( .A(n19881), .B(n19880), .Y(n21541) );
  AOI22XL U24787 ( .A0(n20978), .A1(conv_1[289]), .B0(n22759), .B1(conv_1[274]), .Y(n19882) );
  NAND2XL U24788 ( .A(n19883), .B(n19882), .Y(n21547) );
  AOI22XL U24789 ( .A0(n28528), .A1(n21541), .B0(n34961), .B1(n21547), .Y(
        n19889) );
  AOI22XL U24790 ( .A0(n20978), .A1(conv_1[169]), .B0(n16673), .B1(conv_1[199]), .Y(n19885) );
  NAND2XL U24791 ( .A(n19885), .B(n19884), .Y(n21545) );
  AOI22XL U24792 ( .A0(n20978), .A1(conv_1[349]), .B0(n16673), .B1(conv_1[379]), .Y(n19887) );
  AOI22XL U24793 ( .A0(n16662), .A1(conv_1[364]), .B0(n22690), .B1(conv_1[334]), .Y(n19886) );
  NAND2XL U24794 ( .A(n19887), .B(n19886), .Y(n21546) );
  AOI22XL U24795 ( .A0(n16667), .A1(n21545), .B0(n35234), .B1(n21546), .Y(
        n19888) );
  NAND4XL U24796 ( .A(n19891), .B(n19890), .C(n19889), .D(n19888), .Y(n19892)
         );
  AOI211XL U24797 ( .A0(n28465), .A1(n20245), .B0(n19893), .C0(n19892), .Y(
        n20162) );
  INVXL U24798 ( .A(conv_1[504]), .Y(n27124) );
  INVXL U24799 ( .A(conv_1[489]), .Y(n29987) );
  AOI22XL U24800 ( .A0(n20735), .A1(n27124), .B0(n29987), .B1(n19253), .Y(
        n22521) );
  INVXL U24801 ( .A(conv_1[534]), .Y(n29220) );
  INVXL U24802 ( .A(conv_1[519]), .Y(n30264) );
  AOI22XL U24803 ( .A0(n20735), .A1(n29220), .B0(n30264), .B1(n19253), .Y(
        n22522) );
  AOI22XL U24804 ( .A0(n34950), .A1(n22521), .B0(n21998), .B1(n22522), .Y(
        n19911) );
  INVXL U24805 ( .A(conv_1[264]), .Y(n29201) );
  INVXL U24806 ( .A(conv_1[249]), .Y(n23840) );
  AOI22XL U24807 ( .A0(n20735), .A1(n29201), .B0(n23840), .B1(n19253), .Y(
        n22525) );
  AOI22XL U24808 ( .A0(n22011), .A1(n22525), .B0(n34952), .B1(n22532), .Y(
        n19910) );
  INVXL U24809 ( .A(conv_1[69]), .Y(n27099) );
  INVXL U24810 ( .A(conv_1[54]), .Y(n35311) );
  INVXL U24811 ( .A(conv_1[39]), .Y(n27311) );
  OAI22XL U24812 ( .A0(n22546), .A1(n35311), .B0(n22717), .B1(n27311), .Y(
        n19894) );
  AOI211XL U24813 ( .A0(conv_1[84]), .A1(n16673), .B0(n19895), .C0(n19894), 
        .Y(n21659) );
  INVXL U24814 ( .A(conv_1[159]), .Y(n23398) );
  INVXL U24815 ( .A(conv_1[189]), .Y(n25064) );
  INVXL U24816 ( .A(conv_1[204]), .Y(n31112) );
  OAI22XL U24817 ( .A0(n22612), .A1(n25064), .B0(n24039), .B1(n31112), .Y(
        n19896) );
  AOI211XL U24818 ( .A0(conv_1[174]), .A1(n21011), .B0(n19897), .C0(n19896), 
        .Y(n21664) );
  OAI22XL U24819 ( .A0(n21659), .A1(n28575), .B0(n21664), .B1(n28577), .Y(
        n19908) );
  INVXL U24820 ( .A(conv_1[99]), .Y(n26796) );
  INVXL U24821 ( .A(conv_1[114]), .Y(n31348) );
  INVXL U24822 ( .A(conv_1[129]), .Y(n26714) );
  OAI22XL U24823 ( .A0(n22546), .A1(n31348), .B0(n22612), .B1(n26714), .Y(
        n19898) );
  AOI211XL U24824 ( .A0(conv_1[144]), .A1(n16723), .B0(n19899), .C0(n19898), 
        .Y(n21663) );
  OAI22XL U24825 ( .A0(n21663), .A1(n28479), .B0(n19767), .B1(n21657), .Y(
        n19907) );
  INVXL U24826 ( .A(conv_1[219]), .Y(n34543) );
  INVXL U24827 ( .A(conv_1[234]), .Y(n35407) );
  OAI22XL U24828 ( .A0(n34543), .A1(n22030), .B0(n35407), .B1(n22008), .Y(
        n19906) );
  INVXL U24829 ( .A(conv_1[354]), .Y(n35444) );
  INVXL U24830 ( .A(conv_1[369]), .Y(n23150) );
  OAI22XL U24831 ( .A0(n22546), .A1(n35444), .B0(n22612), .B1(n23150), .Y(
        n19901) );
  INVXL U24832 ( .A(conv_1[339]), .Y(n23015) );
  OAI22XL U24833 ( .A0(n16668), .A1(n23015), .B0(n24039), .B1(n34340), .Y(
        n19900) );
  INVXL U24834 ( .A(conv_1[294]), .Y(n23186) );
  INVXL U24835 ( .A(conv_1[309]), .Y(n24167) );
  INVXL U24836 ( .A(conv_1[324]), .Y(n23314) );
  OAI22XL U24837 ( .A0(n22612), .A1(n24167), .B0(n24039), .B1(n23314), .Y(
        n19903) );
  AOI211XL U24838 ( .A0(conv_1[279]), .A1(n22759), .B0(n19904), .C0(n19903), 
        .Y(n21660) );
  OAI22XL U24839 ( .A0(n21662), .A1(n35196), .B0(n21660), .B1(n18196), .Y(
        n19905) );
  NOR4XL U24840 ( .A(n19908), .B(n19907), .C(n19906), .D(n19905), .Y(n19909)
         );
  NAND3XL U24841 ( .A(n19911), .B(n19910), .C(n19909), .Y(n20087) );
  AOI22XL U24842 ( .A0(n20735), .A1(conv_1[505]), .B0(conv_1[490]), .B1(n18526), .Y(n22488) );
  AOI22XL U24843 ( .A0(n20735), .A1(conv_1[535]), .B0(conv_1[520]), .B1(n18634), .Y(n22489) );
  OAI22XL U24844 ( .A0(n22488), .A1(n21960), .B0(n22489), .B1(n21959), .Y(
        n19929) );
  AOI22XL U24845 ( .A0(n20978), .A1(conv_1[55]), .B0(n16673), .B1(conv_1[85]), 
        .Y(n19913) );
  AOI22XL U24846 ( .A0(n16662), .A1(conv_1[70]), .B0(n22759), .B1(conv_1[40]), 
        .Y(n19912) );
  NAND2XL U24847 ( .A(n19913), .B(n19912), .Y(n21644) );
  INVXL U24848 ( .A(conv_1[370]), .Y(n23155) );
  INVXL U24849 ( .A(conv_1[355]), .Y(n28808) );
  INVXL U24850 ( .A(conv_1[340]), .Y(n23009) );
  OAI22XL U24851 ( .A0(n19902), .A1(n28808), .B0(n22717), .B1(n23009), .Y(
        n19914) );
  AOI211XL U24852 ( .A0(conv_1[385]), .A1(n16673), .B0(n19915), .C0(n19914), 
        .Y(n21637) );
  INVXL U24853 ( .A(conv_1[265]), .Y(n30194) );
  INVXL U24854 ( .A(conv_1[250]), .Y(n35416) );
  AOI22XL U24855 ( .A0(n20735), .A1(n30194), .B0(n35416), .B1(n18634), .Y(
        n22487) );
  AOI22XL U24856 ( .A0(conv_1[235]), .A1(n21999), .B0(n22011), .B1(n22487), 
        .Y(n19927) );
  AOI22XL U24857 ( .A0(n25289), .A1(conv_1[310]), .B0(n16673), .B1(conv_1[325]), .Y(n19917) );
  AOI22XL U24858 ( .A0(n20978), .A1(conv_1[295]), .B0(n25299), .B1(conv_1[280]), .Y(n19916) );
  NAND2XL U24859 ( .A(n19917), .B(n19916), .Y(n21651) );
  INVXL U24860 ( .A(conv_1[115]), .Y(n34561) );
  INVXL U24861 ( .A(conv_1[100]), .Y(n26801) );
  OAI22XL U24862 ( .A0(n22546), .A1(n34561), .B0(n16668), .B1(n26801), .Y(
        n19919) );
  OAI22XL U24863 ( .A0(n21642), .A1(n19767), .B0(n21636), .B1(n28479), .Y(
        n19925) );
  INVXL U24864 ( .A(conv_1[205]), .Y(n35381) );
  INVXL U24865 ( .A(conv_1[190]), .Y(n35367) );
  INVXL U24866 ( .A(conv_1[160]), .Y(n23392) );
  OAI22XL U24867 ( .A0(n22612), .A1(n35367), .B0(n22550), .B1(n23392), .Y(
        n19921) );
  AOI22XL U24868 ( .A0(conv_1[220]), .A1(n16744), .B0(n34952), .B1(n22490), 
        .Y(n19923) );
  OAI21XL U24869 ( .A0(n21654), .A1(n28577), .B0(n19923), .Y(n19924) );
  AOI211XL U24870 ( .A0(n34961), .A1(n21651), .B0(n19925), .C0(n19924), .Y(
        n19926) );
  NAND4BXL U24871 ( .AN(n19929), .B(n19928), .C(n19927), .D(n19926), .Y(n20088) );
  INVXL U24872 ( .A(conv_1[471]), .Y(n27183) );
  INVXL U24873 ( .A(conv_1[456]), .Y(n30023) );
  AOI22XL U24874 ( .A0(n20735), .A1(n27183), .B0(n30023), .B1(n19253), .Y(
        n22460) );
  AOI22XL U24875 ( .A0(n21990), .A1(conv_1[426]), .B0(n21991), .B1(n22460), 
        .Y(n19933) );
  AOI22XL U24876 ( .A0(n21887), .A1(conv_1[441]), .B0(n21954), .B1(conv_1[396]), .Y(n19932) );
  AOI22XL U24877 ( .A0(conv_1[21]), .A1(n22015), .B0(n16734), .B1(conv_1[411]), 
        .Y(n19931) );
  NAND2XL U24878 ( .A(conv_1[6]), .B(n21992), .Y(n19930) );
  NAND4XL U24879 ( .A(n19933), .B(n19932), .C(n19931), .D(n19930), .Y(n20250)
         );
  NAND2XL U24880 ( .A(n22713), .B(n22460), .Y(n20246) );
  INVXL U24881 ( .A(conv_1[531]), .Y(n29244) );
  INVXL U24882 ( .A(conv_1[516]), .Y(n27271) );
  AOI22XL U24883 ( .A0(n20735), .A1(n29244), .B0(n27271), .B1(n19253), .Y(
        n22464) );
  INVXL U24884 ( .A(conv_1[261]), .Y(n29207) );
  INVXL U24885 ( .A(conv_1[246]), .Y(n34333) );
  AOI22XL U24886 ( .A0(n20735), .A1(n29207), .B0(n34333), .B1(n19253), .Y(
        n22471) );
  AOI22XL U24887 ( .A0(n21998), .A1(n22464), .B0(n22011), .B1(n22471), .Y(
        n19934) );
  OAI21XL U24888 ( .A0(n26274), .A1(n20246), .B0(n19934), .Y(n19950) );
  INVXL U24889 ( .A(conv_1[366]), .Y(n22816) );
  INVXL U24890 ( .A(conv_1[336]), .Y(n22987) );
  INVXL U24891 ( .A(conv_1[381]), .Y(n23139) );
  OAI22XL U24892 ( .A0(n22717), .A1(n22987), .B0(n24039), .B1(n23139), .Y(
        n19935) );
  AOI211XL U24893 ( .A0(conv_1[351]), .A1(n25306), .B0(n19936), .C0(n19935), 
        .Y(n21561) );
  INVXL U24894 ( .A(conv_1[51]), .Y(n27315) );
  INVXL U24895 ( .A(conv_1[36]), .Y(n35284) );
  OAI22XL U24896 ( .A0(n22546), .A1(n27315), .B0(n22550), .B1(n35284), .Y(
        n19938) );
  INVXL U24897 ( .A(conv_1[66]), .Y(n27105) );
  INVXL U24898 ( .A(conv_1[81]), .Y(n22871) );
  OAI22XL U24899 ( .A0(n22612), .A1(n27105), .B0(n24039), .B1(n22871), .Y(
        n19937) );
  OAI22XL U24900 ( .A0(n21561), .A1(n35196), .B0(n21560), .B1(n28575), .Y(
        n19948) );
  INVXL U24901 ( .A(conv_1[501]), .Y(n26339) );
  INVXL U24902 ( .A(conv_1[486]), .Y(n35529) );
  AOI22XL U24903 ( .A0(n20735), .A1(n26339), .B0(n35529), .B1(n18526), .Y(
        n22463) );
  AOI22XL U24904 ( .A0(conv_1[231]), .A1(n21999), .B0(n34950), .B1(n22463), 
        .Y(n19947) );
  AOI22XL U24905 ( .A0(n20978), .A1(conv_1[111]), .B0(n22616), .B1(conv_1[96]), 
        .Y(n19940) );
  NAND2XL U24906 ( .A(n19940), .B(n19939), .Y(n21563) );
  AOI22XL U24907 ( .A0(n20978), .A1(conv_1[171]), .B0(n16662), .B1(conv_1[186]), .Y(n19941) );
  NAND2XL U24908 ( .A(n19942), .B(n19941), .Y(n21557) );
  AOI22XL U24909 ( .A0(n28528), .A1(n21563), .B0(n16667), .B1(n21557), .Y(
        n19946) );
  AOI22XL U24910 ( .A0(n20978), .A1(conv_1[291]), .B0(n16662), .B1(conv_1[306]), .Y(n19943) );
  NAND2XL U24911 ( .A(n19944), .B(n19943), .Y(n21562) );
  NAND2XL U24912 ( .A(n22765), .B(n22464), .Y(n21565) );
  NAND2XL U24913 ( .A(n21565), .B(n21566), .Y(n21570) );
  AOI22XL U24914 ( .A0(n34961), .A1(n21562), .B0(n21570), .B1(n24056), .Y(
        n19945) );
  NAND4BXL U24915 ( .AN(n19948), .B(n19947), .C(n19946), .D(n19945), .Y(n19949) );
  AOI211XL U24916 ( .A0(conv_1[216]), .A1(n16744), .B0(n19950), .C0(n19949), 
        .Y(n19951) );
  OAI2BB1XL U24917 ( .A0N(n16700), .A1N(n20250), .B0(n19951), .Y(n20036) );
  NAND2XL U24918 ( .A(n19953), .B(n19952), .Y(n21679) );
  INVXL U24919 ( .A(conv_1[506]), .Y(n27113) );
  INVXL U24920 ( .A(conv_1[491]), .Y(n33208) );
  AOI22XL U24921 ( .A0(n20735), .A1(n27113), .B0(n33208), .B1(n18516), .Y(
        n22595) );
  OAI22XL U24922 ( .A0(n19253), .A1(conv_1[536]), .B0(conv_1[521]), .B1(n35269), .Y(n21689) );
  INVXL U24923 ( .A(n21689), .Y(n22596) );
  AOI22XL U24924 ( .A0(n34950), .A1(n22595), .B0(n34952), .B1(n22590), .Y(
        n19954) );
  OAI21XL U24925 ( .A0(n19767), .A1(n21677), .B0(n19954), .Y(n19968) );
  AOI22XL U24926 ( .A0(n16662), .A1(conv_1[131]), .B0(n22690), .B1(conv_1[101]), .Y(n19955) );
  NAND2XL U24927 ( .A(n19956), .B(n19955), .Y(n21674) );
  NAND2XL U24928 ( .A(n19958), .B(n19957), .Y(n21687) );
  NAND2XL U24929 ( .A(n19960), .B(n19959), .Y(n21686) );
  NAND2XL U24930 ( .A(n19962), .B(n19961), .Y(n21673) );
  AOI22XL U24931 ( .A0(n34961), .A1(n21686), .B0(n35234), .B1(n21673), .Y(
        n19965) );
  AOI22XL U24932 ( .A0(conv_1[221]), .A1(n16744), .B0(n21998), .B1(n22596), 
        .Y(n19964) );
  INVXL U24933 ( .A(conv_1[266]), .Y(n29326) );
  INVXL U24934 ( .A(conv_1[251]), .Y(n26496) );
  AOI22XL U24935 ( .A0(n20735), .A1(n29326), .B0(n26496), .B1(n18526), .Y(
        n22599) );
  AOI22XL U24936 ( .A0(conv_1[236]), .A1(n21999), .B0(n22011), .B1(n22599), 
        .Y(n19963) );
  NAND4XL U24937 ( .A(n19966), .B(n19965), .C(n19964), .D(n19963), .Y(n19967)
         );
  AOI22XL U24938 ( .A0(n20735), .A1(conv_1[503]), .B0(conv_1[488]), .B1(n18634), .Y(n22555) );
  OAI22XL U24939 ( .A0(n18634), .A1(conv_1[263]), .B0(conv_1[248]), .B1(n35269), .Y(n21617) );
  INVXL U24940 ( .A(n21617), .Y(n22557) );
  AOI22XL U24941 ( .A0(n34952), .A1(n22560), .B0(n22011), .B1(n22557), .Y(
        n19969) );
  OAI21XL U24942 ( .A0(n22555), .A1(n21960), .B0(n19969), .Y(n19985) );
  AOI22XL U24943 ( .A0(n16662), .A1(conv_1[128]), .B0(n22690), .B1(conv_1[98]), 
        .Y(n19971) );
  NAND2XL U24944 ( .A(n19971), .B(n19970), .Y(n21625) );
  AOI22XL U24945 ( .A0(n20735), .A1(conv_1[533]), .B0(conv_1[518]), .B1(n18526), .Y(n22556) );
  AOI22XL U24946 ( .A0(n28528), .A1(n21625), .B0(n21623), .B1(n24056), .Y(
        n19983) );
  NAND2XL U24947 ( .A(n19973), .B(n19972), .Y(n21627) );
  AOI22XL U24948 ( .A0(n16662), .A1(conv_1[368]), .B0(n22759), .B1(conv_1[338]), .Y(n19975) );
  NAND2XL U24949 ( .A(n19975), .B(n19974), .Y(n21624) );
  AOI2BB2XL U24950 ( .B0(n21999), .B1(conv_1[233]), .A0N(n21959), .A1N(n22556), 
        .Y(n19981) );
  NAND2XL U24951 ( .A(n19977), .B(n19976), .Y(n21622) );
  NAND2XL U24952 ( .A(n19979), .B(n19978), .Y(n21626) );
  AOI22XL U24953 ( .A0(n16667), .A1(n21622), .B0(n34961), .B1(n21626), .Y(
        n19980) );
  NAND4XL U24954 ( .A(n19983), .B(n19982), .C(n19981), .D(n19980), .Y(n19984)
         );
  AOI211XL U24955 ( .A0(conv_1[218]), .A1(n16744), .B0(n19985), .C0(n19984), 
        .Y(n20041) );
  AOI22XL U24956 ( .A0(n16734), .A1(conv_1[412]), .B0(n21954), .B1(conv_1[397]), .Y(n19989) );
  INVXL U24957 ( .A(conv_1[457]), .Y(n30055) );
  AOI22XL U24958 ( .A0(n20735), .A1(n27604), .B0(n30055), .B1(n18516), .Y(
        n22611) );
  AOI22XL U24959 ( .A0(n21887), .A1(conv_1[442]), .B0(n21991), .B1(n22611), 
        .Y(n19988) );
  AOI22XL U24960 ( .A0(n21990), .A1(conv_1[427]), .B0(conv_1[7]), .B1(n21992), 
        .Y(n19987) );
  NAND2XL U24961 ( .A(conv_1[22]), .B(n22015), .Y(n19986) );
  NAND4XL U24962 ( .A(n19989), .B(n19988), .C(n19987), .D(n19986), .Y(n20272)
         );
  INVXL U24963 ( .A(conv_1[532]), .Y(n29213) );
  INVXL U24964 ( .A(conv_1[517]), .Y(n24917) );
  AOI22XL U24965 ( .A0(n20735), .A1(n29213), .B0(n24917), .B1(n18516), .Y(
        n22627) );
  AOI22XL U24966 ( .A0(n21998), .A1(n22627), .B0(n34952), .B1(n22611), .Y(
        n19991) );
  INVXL U24967 ( .A(conv_1[262]), .Y(n29195) );
  AOI2BB2XL U24968 ( .B0(n20735), .B1(n29195), .A0N(conv_1[247]), .A1N(n35269), 
        .Y(n22623) );
  INVXL U24969 ( .A(n21581), .Y(n20263) );
  AOI22XL U24970 ( .A0(conv_1[232]), .A1(n21999), .B0(n20263), .B1(n34984), 
        .Y(n19990) );
  NAND2XL U24971 ( .A(n19991), .B(n19990), .Y(n20007) );
  INVXL U24972 ( .A(conv_1[487]), .Y(n35536) );
  AOI2BB2XL U24973 ( .B0(n35536), .B1(n18516), .A0N(n18526), .A1N(conv_1[502]), 
        .Y(n22626) );
  AOI22XL U24974 ( .A0(conv_1[217]), .A1(n16744), .B0(n34950), .B1(n22626), 
        .Y(n20005) );
  AOI22XL U24975 ( .A0(n16662), .A1(conv_1[127]), .B0(n22690), .B1(conv_1[97]), 
        .Y(n19992) );
  NAND2XL U24976 ( .A(n19993), .B(n19992), .Y(n21580) );
  AOI22XL U24977 ( .A0(n22759), .A1(conv_1[37]), .B0(n16673), .B1(conv_1[82]), 
        .Y(n19994) );
  NAND2XL U24978 ( .A(n19995), .B(n19994), .Y(n21585) );
  AOI22XL U24979 ( .A0(n16662), .A1(conv_1[187]), .B0(n22690), .B1(conv_1[157]), .Y(n19997) );
  NAND2XL U24980 ( .A(n19997), .B(n19996), .Y(n21597) );
  NAND2XL U24981 ( .A(n22713), .B(n22627), .Y(n21583) );
  OAI2BB1XL U24982 ( .A0N(n36246), .A1N(n22626), .B0(n21583), .Y(n21584) );
  AOI22XL U24983 ( .A0(n16667), .A1(n21597), .B0(n21584), .B1(n24056), .Y(
        n20003) );
  AOI22XL U24984 ( .A0(n16662), .A1(conv_1[307]), .B0(n22690), .B1(conv_1[277]), .Y(n19999) );
  NAND2XL U24985 ( .A(n19999), .B(n19998), .Y(n21579) );
  AOI22XL U24986 ( .A0(n22762), .A1(conv_1[352]), .B0(n16673), .B1(conv_1[382]), .Y(n20001) );
  AOI22XL U24987 ( .A0(n16662), .A1(conv_1[367]), .B0(n22616), .B1(conv_1[337]), .Y(n20000) );
  NAND2XL U24988 ( .A(n20001), .B(n20000), .Y(n21586) );
  AOI22XL U24989 ( .A0(n34961), .A1(n21579), .B0(n35234), .B1(n21586), .Y(
        n20002) );
  NAND4XL U24990 ( .A(n20005), .B(n20004), .C(n20003), .D(n20002), .Y(n20006)
         );
  AOI211XL U24991 ( .A0(n28465), .A1(n20272), .B0(n20007), .C0(n20006), .Y(
        n20035) );
  AOI22XL U24992 ( .A0(n21990), .A1(conv_1[425]), .B0(n21954), .B1(conv_1[395]), .Y(n20012) );
  AOI22XL U24993 ( .A0(n16734), .A1(conv_1[410]), .B0(n21887), .B1(conv_1[440]), .Y(n20011) );
  INVXL U24994 ( .A(conv_1[455]), .Y(n27248) );
  AOI22XL U24995 ( .A0(n20735), .A1(n20008), .B0(n27248), .B1(n18516), .Y(
        n22568) );
  AOI22XL U24996 ( .A0(conv_1[20]), .A1(n22015), .B0(n21991), .B1(n22568), .Y(
        n20010) );
  NAND2XL U24997 ( .A(conv_1[5]), .B(n21992), .Y(n20009) );
  NAND4XL U24998 ( .A(n20012), .B(n20011), .C(n20010), .D(n20009), .Y(n20262)
         );
  AOI22XL U24999 ( .A0(n20735), .A1(conv_1[530]), .B0(conv_1[515]), .B1(n18634), .Y(n22579) );
  INVXL U25000 ( .A(conv_1[260]), .Y(n27561) );
  INVXL U25001 ( .A(conv_1[245]), .Y(n23846) );
  AOI22XL U25002 ( .A0(n20735), .A1(n27561), .B0(n23846), .B1(n18526), .Y(
        n22582) );
  AOI22XL U25003 ( .A0(conv_1[230]), .A1(n21999), .B0(n22011), .B1(n22582), 
        .Y(n20014) );
  NAND2XL U25004 ( .A(n34952), .B(n22568), .Y(n20013) );
  OAI211XL U25005 ( .A0(n22579), .A1(n21959), .B0(n20014), .C0(n20013), .Y(
        n20030) );
  AOI22XL U25006 ( .A0(n20735), .A1(conv_1[500]), .B0(conv_1[485]), .B1(n18526), .Y(n22578) );
  AOI2BB2XL U25007 ( .B0(conv_1[215]), .B1(n16744), .A0N(n21960), .A1N(n22578), 
        .Y(n20028) );
  AOI22XL U25008 ( .A0(n16662), .A1(conv_1[125]), .B0(n22616), .B1(conv_1[95]), 
        .Y(n20016) );
  NAND2XL U25009 ( .A(n20016), .B(n20015), .Y(n21599) );
  AOI22XL U25010 ( .A0(n22762), .A1(conv_1[170]), .B0(n16662), .B1(conv_1[185]), .Y(n20018) );
  AOI22XL U25011 ( .A0(n18658), .A1(conv_1[155]), .B0(n16673), .B1(conv_1[200]), .Y(n20017) );
  NAND2XL U25012 ( .A(n20018), .B(n20017), .Y(n21601) );
  AOI22XL U25013 ( .A0(n28528), .A1(n21599), .B0(n16667), .B1(n21601), .Y(
        n20027) );
  AOI22XL U25014 ( .A0(n22770), .A1(conv_1[50]), .B0(n16673), .B1(conv_1[80]), 
        .Y(n20020) );
  AOI22XL U25015 ( .A0(n16662), .A1(conv_1[65]), .B0(n25299), .B1(conv_1[35]), 
        .Y(n20019) );
  NAND2XL U25016 ( .A(n20020), .B(n20019), .Y(n21610) );
  AOI22XL U25017 ( .A0(n16662), .A1(conv_1[305]), .B0(n22759), .B1(conv_1[275]), .Y(n20022) );
  AOI22XL U25018 ( .A0(n22762), .A1(conv_1[290]), .B0(n16673), .B1(conv_1[320]), .Y(n20021) );
  NAND2XL U25019 ( .A(n20022), .B(n20021), .Y(n21598) );
  AOI22XL U25020 ( .A0(n25299), .A1(conv_1[335]), .B0(n16673), .B1(conv_1[380]), .Y(n20024) );
  AOI22XL U25021 ( .A0(n22770), .A1(conv_1[350]), .B0(n16662), .B1(conv_1[365]), .Y(n20023) );
  NAND2XL U25022 ( .A(n20024), .B(n20023), .Y(n21605) );
  AOI22XL U25023 ( .A0(n34961), .A1(n21598), .B0(n35234), .B1(n21605), .Y(
        n20025) );
  NAND4XL U25024 ( .A(n20028), .B(n20027), .C(n20026), .D(n20025), .Y(n20029)
         );
  AOI211XL U25025 ( .A0(n28465), .A1(n20262), .B0(n20030), .C0(n20029), .Y(
        n20034) );
  NAND4XL U25026 ( .A(n20040), .B(n20041), .C(n20035), .D(n20034), .Y(n20031)
         );
  NOR4XL U25027 ( .A(n20087), .B(n20088), .C(n20036), .D(n20031), .Y(n20032)
         );
  OAI211XL U25028 ( .A0(n20033), .A1(n35135), .B0(n20162), .C0(n20032), .Y(
        n20038) );
  NOR4BBXL U25029 ( .AN(n20087), .BN(n20088), .C(n20040), .D(n20041), .Y(
        n20092) );
  INVXL U25030 ( .A(n20281), .Y(n20042) );
  AOI22XL U25031 ( .A0(n20042), .A1(n20041), .B0(n20287), .B1(n20040), .Y(
        n20091) );
  INVXL U25032 ( .A(conv_1[508]), .Y(n27184) );
  INVXL U25033 ( .A(conv_1[493]), .Y(n33352) );
  AOI22XL U25034 ( .A0(n35269), .A1(n27184), .B0(n33352), .B1(n18634), .Y(
        n22766) );
  AOI22XL U25035 ( .A0(conv_1[238]), .A1(n21999), .B0(n34950), .B1(n22766), 
        .Y(n20056) );
  AOI22XL U25036 ( .A0(n16716), .A1(conv_1[193]), .B0(n16673), .B1(conv_1[208]), .Y(n20044) );
  AOI22XL U25037 ( .A0(n22762), .A1(conv_1[178]), .B0(n22690), .B1(conv_1[163]), .Y(n20043) );
  NAND2XL U25038 ( .A(n20044), .B(n20043), .Y(n21728) );
  AOI22XL U25039 ( .A0(n22616), .A1(conv_1[283]), .B0(n16673), .B1(conv_1[328]), .Y(n20046) );
  AOI22XL U25040 ( .A0(n22762), .A1(conv_1[298]), .B0(n16662), .B1(conv_1[313]), .Y(n20045) );
  NAND2XL U25041 ( .A(n20046), .B(n20045), .Y(n21732) );
  AOI22XL U25042 ( .A0(n16667), .A1(n21728), .B0(n34961), .B1(n21732), .Y(
        n20055) );
  AOI22XL U25043 ( .A0(n25299), .A1(conv_1[103]), .B0(n16673), .B1(conv_1[148]), .Y(n20048) );
  NAND2XL U25044 ( .A(n20048), .B(n20047), .Y(n21734) );
  AOI22XL U25045 ( .A0(n22759), .A1(conv_1[43]), .B0(n16673), .B1(conv_1[88]), 
        .Y(n20049) );
  NAND2XL U25046 ( .A(n20050), .B(n20049), .Y(n21727) );
  AOI22XL U25047 ( .A0(n22770), .A1(conv_1[358]), .B0(n16662), .B1(conv_1[373]), .Y(n20052) );
  AOI22XL U25048 ( .A0(n25299), .A1(conv_1[343]), .B0(n16673), .B1(conv_1[388]), .Y(n20051) );
  NAND2XL U25049 ( .A(n20052), .B(n20051), .Y(n21733) );
  INVXL U25050 ( .A(conv_1[538]), .Y(n27999) );
  INVXL U25051 ( .A(conv_1[523]), .Y(n30261) );
  AOI22XL U25052 ( .A0(n35269), .A1(n27999), .B0(n30261), .B1(n18516), .Y(
        n22767) );
  NAND2XL U25053 ( .A(n22713), .B(n22767), .Y(n20333) );
  NAND2XL U25054 ( .A(n20333), .B(n21726), .Y(n21735) );
  AOI22XL U25055 ( .A0(n35234), .A1(n21733), .B0(n21735), .B1(n24056), .Y(
        n20053) );
  NAND4XL U25056 ( .A(n20056), .B(n20055), .C(n20054), .D(n20053), .Y(n20064)
         );
  INVXL U25057 ( .A(conv_1[28]), .Y(n33436) );
  INVXL U25058 ( .A(conv_1[13]), .Y(n27362) );
  INVXL U25059 ( .A(conv_1[478]), .Y(n33248) );
  INVXL U25060 ( .A(conv_1[463]), .Y(n28747) );
  AOI22XL U25061 ( .A0(n35269), .A1(n33248), .B0(n28747), .B1(n18526), .Y(
        n22771) );
  AOI22XL U25062 ( .A0(n21990), .A1(conv_1[433]), .B0(n21991), .B1(n22771), 
        .Y(n20058) );
  AOI22XL U25063 ( .A0(n16734), .A1(conv_1[418]), .B0(n21954), .B1(conv_1[403]), .Y(n20057) );
  OAI211XL U25064 ( .A0(n27362), .A1(n22018), .B0(n20058), .C0(n20057), .Y(
        n20059) );
  AOI211XL U25065 ( .A0(conv_1[448]), .A1(n21887), .B0(n20060), .C0(n20059), 
        .Y(n20336) );
  INVXL U25066 ( .A(conv_1[268]), .Y(n34083) );
  INVXL U25067 ( .A(conv_1[253]), .Y(n27981) );
  AOI22XL U25068 ( .A0(n35269), .A1(n34083), .B0(n27981), .B1(n18634), .Y(
        n22772) );
  AOI22XL U25069 ( .A0(n22011), .A1(n22772), .B0(n21998), .B1(n22767), .Y(
        n20062) );
  AOI22XL U25070 ( .A0(conv_1[223]), .A1(n16744), .B0(n34952), .B1(n22771), 
        .Y(n20061) );
  OAI211XL U25071 ( .A0(n20336), .A1(n35135), .B0(n20062), .C0(n20061), .Y(
        n20063) );
  AOI22XL U25072 ( .A0(n21990), .A1(conv_1[432]), .B0(n21887), .B1(conv_1[447]), .Y(n20068) );
  INVXL U25073 ( .A(conv_1[477]), .Y(n29828) );
  INVXL U25074 ( .A(conv_1[462]), .Y(n28730) );
  AOI22XL U25075 ( .A0(n20735), .A1(n29828), .B0(n28730), .B1(n18634), .Y(
        n22732) );
  AOI22XL U25076 ( .A0(n21954), .A1(conv_1[402]), .B0(n21991), .B1(n22732), 
        .Y(n20067) );
  AOI22XL U25077 ( .A0(conv_1[27]), .A1(n22015), .B0(n16734), .B1(conv_1[417]), 
        .Y(n20066) );
  NAND2XL U25078 ( .A(conv_1[12]), .B(n21992), .Y(n20065) );
  NAND4XL U25079 ( .A(n20068), .B(n20067), .C(n20066), .D(n20065), .Y(n20327)
         );
  AOI22XL U25080 ( .A0(n35269), .A1(conv_1[537]), .B0(conv_1[522]), .B1(n18634), .Y(n22745) );
  AOI22XL U25081 ( .A0(n35269), .A1(conv_1[507]), .B0(conv_1[492]), .B1(n19253), .Y(n22744) );
  AOI22XL U25082 ( .A0(n35236), .A1(n21768), .B0(n34952), .B1(n22732), .Y(
        n20072) );
  AOI22XL U25083 ( .A0(n22762), .A1(conv_1[357]), .B0(n16662), .B1(conv_1[372]), .Y(n20070) );
  AOI22XL U25084 ( .A0(n22616), .A1(conv_1[342]), .B0(n16673), .B1(conv_1[387]), .Y(n20069) );
  NAND2XL U25085 ( .A(n20070), .B(n20069), .Y(n21755) );
  NAND2XL U25086 ( .A(n35234), .B(n21755), .Y(n20071) );
  OAI211XL U25087 ( .A0(n21760), .A1(n19767), .B0(n20072), .C0(n20071), .Y(
        n20086) );
  INVXL U25088 ( .A(conv_1[267]), .Y(n29355) );
  INVXL U25089 ( .A(conv_1[252]), .Y(n33665) );
  AOI22XL U25090 ( .A0(n20735), .A1(n29355), .B0(n33665), .B1(n19253), .Y(
        n22735) );
  AOI22XL U25091 ( .A0(conv_1[237]), .A1(n21999), .B0(n22011), .B1(n22735), 
        .Y(n20084) );
  INVXL U25092 ( .A(n22744), .Y(n21750) );
  AOI22XL U25093 ( .A0(conv_1[222]), .A1(n16744), .B0(n34950), .B1(n21750), 
        .Y(n20083) );
  AOI22XL U25094 ( .A0(n16666), .A1(conv_1[177]), .B0(n22690), .B1(conv_1[162]), .Y(n20074) );
  AOI22XL U25095 ( .A0(n16716), .A1(conv_1[192]), .B0(n16673), .B1(conv_1[207]), .Y(n20073) );
  NAND2XL U25096 ( .A(n20074), .B(n20073), .Y(n21775) );
  AOI22XL U25097 ( .A0(n22762), .A1(conv_1[297]), .B0(n18658), .B1(conv_1[282]), .Y(n20076) );
  AOI22XL U25098 ( .A0(n16716), .A1(conv_1[312]), .B0(n16673), .B1(conv_1[327]), .Y(n20075) );
  NAND2XL U25099 ( .A(n20076), .B(n20075), .Y(n21767) );
  AOI22XL U25100 ( .A0(n16667), .A1(n21775), .B0(n34961), .B1(n21767), .Y(
        n20082) );
  AOI22XL U25101 ( .A0(n22762), .A1(conv_1[117]), .B0(n22759), .B1(conv_1[102]), .Y(n20078) );
  AOI22XL U25102 ( .A0(n16716), .A1(conv_1[132]), .B0(n16673), .B1(conv_1[147]), .Y(n20077) );
  NAND2XL U25103 ( .A(n20078), .B(n20077), .Y(n21757) );
  AOI22XL U25104 ( .A0(n25299), .A1(conv_1[42]), .B0(n16673), .B1(conv_1[87]), 
        .Y(n20080) );
  AOI22XL U25105 ( .A0(n22762), .A1(conv_1[57]), .B0(n16662), .B1(conv_1[72]), 
        .Y(n20079) );
  NAND2XL U25106 ( .A(n20080), .B(n20079), .Y(n21754) );
  NAND4XL U25107 ( .A(n20084), .B(n20083), .C(n20082), .D(n20081), .Y(n20085)
         );
  AOI211XL U25108 ( .A0(n28465), .A1(n20327), .B0(n20086), .C0(n20085), .Y(
        n20094) );
  OAI22XL U25109 ( .A0(n20297), .A1(n20088), .B0(n20306), .B1(n20087), .Y(
        n20089) );
  NOR4XL U25110 ( .A(n20093), .B(n20094), .C(n20161), .D(n20089), .Y(n20090)
         );
  OAI211XL U25111 ( .A0(n28465), .A1(n20092), .B0(n20091), .C0(n20090), .Y(
        n20096) );
  AND3XL U25112 ( .A(n20161), .B(n20094), .C(n20093), .Y(n20095) );
  NAND2XL U25113 ( .A(n34800), .B(pool[5]), .Y(n20100) );
  OAI21XL U25114 ( .A0(n20101), .A1(n34800), .B0(n20100), .Y(N29221) );
  ADDFX1 U25115 ( .A(DP_OP_5170J1_126_4278_n64), .B(n20103), .CI(n20102), .CO(
        n20106), .S(n19633) );
  AOI22XL U25116 ( .A0(affine_2[21]), .A1(n33367), .B0(n16674), .B1(n20104), 
        .Y(n20105) );
  NAND2XL U25117 ( .A(n20105), .B(n33350), .Y(n16540) );
  ADDFX1 U25118 ( .A(DP_OP_5170J1_126_4278_n59), .B(DP_OP_5170J1_126_4278_n63), 
        .CI(n20106), .CO(n20112), .S(n20104) );
  AOI22XL U25119 ( .A0(affine_2[24]), .A1(n33367), .B0(n16674), .B1(n20107), 
        .Y(n20108) );
  NAND2XL U25120 ( .A(n20108), .B(n33350), .Y(n16537) );
  ADDFX1 U25121 ( .A(DP_OP_5170J1_126_4278_n44), .B(DP_OP_5170J1_126_4278_n48), 
        .CI(n20109), .CO(n20135), .S(n20107) );
  AOI22XL U25122 ( .A0(affine_2[26]), .A1(n33367), .B0(n16674), .B1(n20110), 
        .Y(n20111) );
  NAND2XL U25123 ( .A(n20111), .B(n33350), .Y(n16535) );
  ADDFX1 U25124 ( .A(DP_OP_5170J1_126_4278_n54), .B(DP_OP_5170J1_126_4278_n58), 
        .CI(n20112), .CO(n20141), .S(n20113) );
  AOI22XL U25125 ( .A0(affine_2[22]), .A1(n33367), .B0(n16674), .B1(n20113), 
        .Y(n20114) );
  NAND2XL U25126 ( .A(n20114), .B(n33350), .Y(n16539) );
  ADDFX1 U25127 ( .A(DP_OP_5171J1_127_4278_n64), .B(n20116), .CI(n20115), .CO(
        n20126), .S(n19713) );
  AOI22XL U25128 ( .A0(affine_2[8]), .A1(n33367), .B0(n16674), .B1(n20117), 
        .Y(n20118) );
  NAND2XL U25129 ( .A(n20118), .B(n33368), .Y(n16571) );
  ADDFX1 U25130 ( .A(DP_OP_5171J1_127_4278_n49), .B(DP_OP_5171J1_127_4278_n53), 
        .CI(n20119), .CO(n20132), .S(n20120) );
  AOI22XL U25131 ( .A0(affine_2[7]), .A1(n33367), .B0(n16674), .B1(n20120), 
        .Y(n20121) );
  NAND2XL U25132 ( .A(n20121), .B(n33368), .Y(n16572) );
  ADDFX1 U25133 ( .A(DP_OP_5169J1_125_4278_n64), .B(n20123), .CI(n20122), .CO(
        n20129), .S(n19734) );
  AOI22XL U25134 ( .A0(affine_2[39]), .A1(n33367), .B0(n16674), .B1(n20124), 
        .Y(n20125) );
  NAND2XL U25135 ( .A(n20125), .B(n33340), .Y(n16554) );
  ADDFX1 U25136 ( .A(DP_OP_5171J1_127_4278_n59), .B(DP_OP_5171J1_127_4278_n63), 
        .CI(n20126), .CO(n20150), .S(n20127) );
  AOI22XL U25137 ( .A0(affine_2[5]), .A1(n33367), .B0(n16674), .B1(n20127), 
        .Y(n20128) );
  NAND2XL U25138 ( .A(n20128), .B(n33368), .Y(n16574) );
  ADDFX1 U25139 ( .A(DP_OP_5169J1_125_4278_n59), .B(DP_OP_5169J1_125_4278_n63), 
        .CI(n20129), .CO(n20156), .S(n20130) );
  AOI22XL U25140 ( .A0(affine_2[37]), .A1(n33367), .B0(n16674), .B1(n20130), 
        .Y(n20131) );
  NAND2XL U25141 ( .A(n20131), .B(n33340), .Y(n16556) );
  ADDFX1 U25142 ( .A(DP_OP_5171J1_127_4278_n44), .B(DP_OP_5171J1_127_4278_n48), 
        .CI(n20132), .CO(n20138), .S(n20117) );
  AOI22XL U25143 ( .A0(affine_2[9]), .A1(n33367), .B0(n16674), .B1(n20133), 
        .Y(n20134) );
  NAND2XL U25144 ( .A(n20134), .B(n33368), .Y(n16570) );
  ADDFX1 U25145 ( .A(DP_OP_5170J1_126_4278_n39), .B(DP_OP_5170J1_126_4278_n43), 
        .CI(n20135), .CO(n20352), .S(n20136) );
  AOI22XL U25146 ( .A0(affine_2[25]), .A1(n33367), .B0(n16674), .B1(n20136), 
        .Y(n20137) );
  NAND2XL U25147 ( .A(n20137), .B(n33350), .Y(n16536) );
  ADDFX1 U25148 ( .A(DP_OP_5171J1_127_4278_n39), .B(DP_OP_5171J1_127_4278_n43), 
        .CI(n20138), .CO(n20182), .S(n20133) );
  AOI22XL U25149 ( .A0(affine_2[10]), .A1(n33367), .B0(n16674), .B1(n20139), 
        .Y(n20140) );
  NAND2XL U25150 ( .A(n20140), .B(n33368), .Y(n16569) );
  ADDFX1 U25151 ( .A(DP_OP_5170J1_126_4278_n49), .B(DP_OP_5170J1_126_4278_n53), 
        .CI(n20141), .CO(n20109), .S(n20142) );
  AOI22XL U25152 ( .A0(affine_2[23]), .A1(n33367), .B0(n16674), .B1(n20142), 
        .Y(n20143) );
  NAND2XL U25153 ( .A(n20143), .B(n33350), .Y(n16538) );
  AOI22XL U25154 ( .A0(affine_2[41]), .A1(n33367), .B0(n16674), .B1(n20145), 
        .Y(n20146) );
  NAND2XL U25155 ( .A(n20146), .B(n33340), .Y(n16552) );
  AOI22XL U25156 ( .A0(affine_2[42]), .A1(n33367), .B0(n16674), .B1(n20148), 
        .Y(n20149) );
  NAND2XL U25157 ( .A(n20149), .B(n33340), .Y(n16551) );
  ADDFX1 U25158 ( .A(DP_OP_5171J1_127_4278_n54), .B(DP_OP_5171J1_127_4278_n58), 
        .CI(n20150), .CO(n20119), .S(n20151) );
  AOI22XL U25159 ( .A0(affine_2[6]), .A1(n33367), .B0(n16674), .B1(n20151), 
        .Y(n20152) );
  NAND2XL U25160 ( .A(n20152), .B(n33368), .Y(n16573) );
  AOI22XL U25161 ( .A0(affine_2[40]), .A1(n33367), .B0(n16674), .B1(n20154), 
        .Y(n20155) );
  NAND2XL U25162 ( .A(n20155), .B(n33340), .Y(n16553) );
  AOI22XL U25163 ( .A0(affine_2[38]), .A1(n33367), .B0(n16674), .B1(n20157), 
        .Y(n20158) );
  NAND2XL U25164 ( .A(n20158), .B(n33340), .Y(n16555) );
  AOI22XL U25165 ( .A0(n34798), .A1(n20160), .B0(n20159), .B1(n34800), .Y(
        N29224) );
  AOI22XL U25166 ( .A0(n34798), .A1(n20162), .B0(n20161), .B1(n34800), .Y(
        N29225) );
  INVXL U25167 ( .A(n36122), .Y(n20360) );
  INVXL U25168 ( .A(filter_3_bias[4]), .Y(n20169) );
  INVXL U25169 ( .A(filter_2_bias[4]), .Y(n36110) );
  AOI22XL U25170 ( .A0(n36114), .A1(n20169), .B0(n36110), .B1(n20180), .Y(
        n14728) );
  INVXL U25171 ( .A(n20179), .Y(n20166) );
  INVXL U25172 ( .A(filter_3_bias[1]), .Y(n20176) );
  AOI22XL U25173 ( .A0(n36114), .A1(n36139), .B0(n20176), .B1(n20180), .Y(
        n14720) );
  INVXL U25174 ( .A(filter_3_bias[3]), .Y(n20173) );
  INVXL U25175 ( .A(filter_2_bias[3]), .Y(n36111) );
  AOI22XL U25176 ( .A0(n36114), .A1(n20173), .B0(n36111), .B1(n20180), .Y(
        n14725) );
  NAND2XL U25177 ( .A(n20179), .B(in_data[10]), .Y(n20178) );
  INVXL U25178 ( .A(in_data[11]), .Y(n20172) );
  NAND2XL U25179 ( .A(n20170), .B(in_data[12]), .Y(n20174) );
  AOI22XL U25180 ( .A0(n36114), .A1(n36148), .B0(n20169), .B1(n20180), .Y(
        n14729) );
  INVXL U25181 ( .A(n20170), .Y(n20171) );
  AOI22XL U25182 ( .A0(n36114), .A1(n36145), .B0(n20173), .B1(n20180), .Y(
        n14726) );
  INVXL U25183 ( .A(filter_3_bias[0]), .Y(n20175) );
  AOI22XL U25184 ( .A0(n36114), .A1(n36124), .B0(n20175), .B1(n20180), .Y(
        n14735) );
  INVXL U25185 ( .A(filter_3_bias[5]), .Y(n20177) );
  AOI22XL U25186 ( .A0(n36114), .A1(n36151), .B0(n20177), .B1(n20180), .Y(
        n14732) );
  INVXL U25187 ( .A(filter_2_bias[0]), .Y(n36108) );
  AOI22XL U25188 ( .A0(n36114), .A1(n20175), .B0(n36108), .B1(n20180), .Y(
        n14734) );
  INVXL U25189 ( .A(filter_2_bias[1]), .Y(n36113) );
  AOI22XL U25190 ( .A0(n36114), .A1(n20176), .B0(n36113), .B1(n20180), .Y(
        n14719) );
  INVXL U25191 ( .A(filter_2_bias[5]), .Y(n36109) );
  AOI22XL U25192 ( .A0(n36114), .A1(n20177), .B0(n36109), .B1(n20180), .Y(
        n14731) );
  INVXL U25193 ( .A(filter_3_bias[2]), .Y(n20181) );
  INVXL U25194 ( .A(filter_2_bias[2]), .Y(n36112) );
  AOI22XL U25195 ( .A0(n36114), .A1(n20181), .B0(n36112), .B1(n20180), .Y(
        n14722) );
  AOI22XL U25196 ( .A0(n36114), .A1(n36142), .B0(n20181), .B1(n20180), .Y(
        n14723) );
  ADDFX1 U25197 ( .A(DP_OP_5171J1_127_4278_n34), .B(DP_OP_5171J1_127_4278_n38), 
        .CI(n20182), .CO(n22092), .S(n20139) );
  AOI22XL U25198 ( .A0(affine_2[11]), .A1(n33367), .B0(n16674), .B1(n20183), 
        .Y(n20184) );
  NAND2XL U25199 ( .A(n20184), .B(n33368), .Y(n16568) );
  AOI22XL U25200 ( .A0(n35236), .A1(n21469), .B0(n16671), .B1(n21459), .Y(
        n20187) );
  OAI211XL U25201 ( .A0(n21466), .A1(n16672), .B0(n20187), .C0(n20186), .Y(
        n20192) );
  AOI22XL U25202 ( .A0(n35195), .A1(n21467), .B0(n34906), .B1(n21468), .Y(
        n20189) );
  AOI22XL U25203 ( .A0(n16660), .A1(n21460), .B0(n19179), .B1(n21458), .Y(
        n20188) );
  OAI211XL U25204 ( .A0(n20190), .A1(n25853), .B0(n20189), .C0(n20188), .Y(
        n20191) );
  INVXL U25205 ( .A(conv_1[239]), .Y(n33852) );
  OAI22XL U25206 ( .A0(n22712), .A1(n25872), .B0(n33852), .B1(n26085), .Y(
        n20198) );
  AOI22XL U25207 ( .A0(n16671), .A1(n21707), .B0(n21708), .B1(n35231), .Y(
        n20196) );
  OAI211XL U25208 ( .A0(n21724), .A1(n35239), .B0(n20196), .C0(n20195), .Y(
        n20197) );
  AOI211XL U25209 ( .A0(n35236), .A1(n21709), .B0(n20198), .C0(n20197), .Y(
        n20203) );
  OAI22XL U25210 ( .A0(n22721), .A1(n26026), .B0(n28606), .B1(n26029), .Y(
        n20200) );
  OAI22XL U25211 ( .A0(n21713), .A1(n35198), .B0(n21705), .B1(n26039), .Y(
        n20199) );
  AOI211XL U25212 ( .A0(n16755), .A1(n20201), .B0(n20200), .C0(n20199), .Y(
        n20202) );
  NAND2XL U25213 ( .A(n20203), .B(n20202), .Y(n20348) );
  AOI22XL U25214 ( .A0(n34903), .A1(n22635), .B0(n26081), .B1(n22638), .Y(
        n20205) );
  NAND2XL U25215 ( .A(conv_1[213]), .B(n26082), .Y(n20204) );
  OAI211XL U25216 ( .A0(n28479), .A1(n20206), .B0(n20205), .C0(n20204), .Y(
        n20213) );
  AOI22XL U25217 ( .A0(conv_1[228]), .A1(n26059), .B0(n26276), .B1(n21479), 
        .Y(n20211) );
  AOI22XL U25218 ( .A0(n19179), .A1(n21481), .B0(n16671), .B1(n21484), .Y(
        n20210) );
  AOI22XL U25219 ( .A0(n16660), .A1(n21483), .B0(n35231), .B1(n21485), .Y(
        n20209) );
  AOI22XL U25220 ( .A0(n35195), .A1(n21480), .B0(n35236), .B1(n21482), .Y(
        n20208) );
  NAND4XL U25221 ( .A(n20211), .B(n20210), .C(n20209), .D(n20208), .Y(n20212)
         );
  OR2XL U25222 ( .A(n22682), .B(n21688), .Y(n21498) );
  AOI22XL U25223 ( .A0(n16671), .A1(n21506), .B0(n35231), .B1(n21501), .Y(
        n20215) );
  AOI32XL U25224 ( .A0(n21498), .A1(n20215), .A2(n21496), .B0(n28479), .B1(
        n20215), .Y(n20222) );
  AOI22XL U25225 ( .A0(conv_1[226]), .A1(n26059), .B0(n26081), .B1(n22696), 
        .Y(n20220) );
  OAI2BB2XL U25226 ( .B0(n22683), .B1(n26026), .A0N(n26082), .A1N(conv_1[211]), 
        .Y(n20217) );
  OAI22XL U25227 ( .A0(n21504), .A1(n35198), .B0(n21503), .B1(n18208), .Y(
        n20216) );
  AOI211XL U25228 ( .A0(n16755), .A1(n20218), .B0(n20217), .C0(n20216), .Y(
        n20219) );
  OAI211XL U25229 ( .A0(n21497), .A1(n35239), .B0(n20220), .C0(n20219), .Y(
        n20221) );
  AOI211XL U25230 ( .A0(n19179), .A1(n21505), .B0(n20222), .C0(n20221), .Y(
        n34841) );
  AOI222XL U25231 ( .A0(n20351), .A1(pool[36]), .B0(n20351), .B1(n34841), .C0(
        pool[36]), .C1(n34841), .Y(n20235) );
  AOI22XL U25232 ( .A0(n35236), .A1(n21519), .B0(conv_1[212]), .B1(n26082), 
        .Y(n20234) );
  AOI22XL U25233 ( .A0(n35195), .A1(n21516), .B0(n16671), .B1(n21521), .Y(
        n20233) );
  OAI22XL U25234 ( .A0(n34989), .A1(n20224), .B0(n25853), .B1(n20223), .Y(
        n20229) );
  AOI22XL U25235 ( .A0(n16659), .A1(n21517), .B0(n34903), .B1(n22662), .Y(
        n20226) );
  AOI22XL U25236 ( .A0(n16660), .A1(n21522), .B0(n19179), .B1(n21515), .Y(
        n20225) );
  OAI211XL U25237 ( .A0(n20227), .A1(n23053), .B0(n20226), .C0(n20225), .Y(
        n20228) );
  AOI211XL U25238 ( .A0(conv_1[227]), .A1(n26059), .B0(n20229), .C0(n20228), 
        .Y(n20232) );
  NAND2XL U25239 ( .A(n16755), .B(n20230), .Y(n20231) );
  AOI222XL U25240 ( .A0(n20235), .A1(n34842), .B0(n20235), .B1(n34843), .C0(
        n34842), .C1(n34843), .Y(n20236) );
  AOI222XL U25241 ( .A0(pool[38]), .A1(n20611), .B0(pool[38]), .B1(n20236), 
        .C0(n20611), .C1(n20236), .Y(n20317) );
  AOI22XL U25242 ( .A0(conv_1[214]), .A1(n26082), .B0(n35231), .B1(n21544), 
        .Y(n20237) );
  OAI21XL U25243 ( .A0(n22498), .A1(n25872), .B0(n20237), .Y(n20244) );
  AOI22XL U25244 ( .A0(conv_1[229]), .A1(n26059), .B0(n25875), .B1(n22510), 
        .Y(n20242) );
  AOI22XL U25245 ( .A0(n35195), .A1(n21543), .B0(n35236), .B1(n21541), .Y(
        n20241) );
  NAND2XL U25246 ( .A(n22765), .B(n22499), .Y(n21537) );
  NAND2XL U25247 ( .A(n21535), .B(n21537), .Y(n20238) );
  AOI22XL U25248 ( .A0(n16659), .A1(n20238), .B0(n16671), .B1(n21547), .Y(
        n20240) );
  AOI22XL U25249 ( .A0(n16660), .A1(n21545), .B0(n19179), .B1(n21546), .Y(
        n20239) );
  NAND4XL U25250 ( .A(n20242), .B(n20241), .C(n20240), .D(n20239), .Y(n20243)
         );
  AOI211XL U25251 ( .A0(n16755), .A1(n20245), .B0(n20244), .C0(n20243), .Y(
        n20609) );
  AOI22XL U25252 ( .A0(n16660), .A1(n21557), .B0(n35231), .B1(n21570), .Y(
        n20247) );
  AOI32XL U25253 ( .A0(n21566), .A1(n20247), .A2(n20246), .B0(n28479), .B1(
        n20247), .Y(n20254) );
  AOI22XL U25254 ( .A0(conv_1[216]), .A1(n26082), .B0(n16671), .B1(n21562), 
        .Y(n20252) );
  INVXL U25255 ( .A(conv_1[231]), .Y(n29267) );
  OAI22XL U25256 ( .A0(n29267), .A1(n26085), .B0(n35196), .B1(n21564), .Y(
        n20249) );
  OAI22XL U25257 ( .A0(n21561), .A1(n26039), .B0(n21560), .B1(n35239), .Y(
        n20248) );
  AOI211XL U25258 ( .A0(n16755), .A1(n20250), .B0(n20249), .C0(n20248), .Y(
        n20251) );
  OAI211XL U25259 ( .A0(n26162), .A1(n21565), .B0(n20252), .C0(n20251), .Y(
        n20253) );
  AOI211XL U25260 ( .A0(n35236), .A1(n21563), .B0(n20254), .C0(n20253), .Y(
        n20273) );
  AOI22XL U25261 ( .A0(n16660), .A1(n21601), .B0(n26081), .B1(n22582), .Y(
        n20255) );
  OAI21XL U25262 ( .A0(n22579), .A1(n26026), .B0(n20255), .Y(n20261) );
  AOI22XL U25263 ( .A0(conv_1[215]), .A1(n26082), .B0(conv_1[230]), .B1(n26059), .Y(n20259) );
  AOI22XL U25264 ( .A0(n21600), .A1(n25879), .B0(n34903), .B1(n22568), .Y(
        n20258) );
  AOI22XL U25265 ( .A0(n19179), .A1(n21605), .B0(n16671), .B1(n21598), .Y(
        n20257) );
  AOI22XL U25266 ( .A0(n35195), .A1(n21610), .B0(n35236), .B1(n21599), .Y(
        n20256) );
  NAND4XL U25267 ( .A(n20259), .B(n20258), .C(n20257), .D(n20256), .Y(n20260)
         );
  AOI211XL U25268 ( .A0(n16755), .A1(n20262), .B0(n20261), .C0(n20260), .Y(
        n20314) );
  AOI22XL U25269 ( .A0(conv_1[232]), .A1(n26059), .B0(n35234), .B1(n20263), 
        .Y(n20265) );
  NAND2XL U25270 ( .A(n26066), .B(n22626), .Y(n20264) );
  OAI211XL U25271 ( .A0(n21583), .A1(n26162), .B0(n20265), .C0(n20264), .Y(
        n20271) );
  AOI22XL U25272 ( .A0(conv_1[217]), .A1(n26082), .B0(n34903), .B1(n22611), 
        .Y(n20269) );
  AOI22XL U25273 ( .A0(n35195), .A1(n21585), .B0(n35231), .B1(n21584), .Y(
        n20268) );
  AOI22XL U25274 ( .A0(n35236), .A1(n21580), .B0(n19179), .B1(n21586), .Y(
        n20267) );
  AOI22XL U25275 ( .A0(n16660), .A1(n21597), .B0(n16671), .B1(n21579), .Y(
        n20266) );
  NAND4XL U25276 ( .A(n20269), .B(n20268), .C(n20267), .D(n20266), .Y(n20270)
         );
  AOI211XL U25277 ( .A0(n16755), .A1(n20272), .B0(n20271), .C0(n20270), .Y(
        n20313) );
  NOR4XL U25278 ( .A(n20609), .B(n20273), .C(n20314), .D(n20313), .Y(n20316)
         );
  AND2XL U25279 ( .A(n20609), .B(n20273), .Y(n20312) );
  AOI22XL U25280 ( .A0(n35236), .A1(n21625), .B0(n26081), .B1(n22557), .Y(
        n20283) );
  INVXL U25281 ( .A(conv_1[218]), .Y(n24684) );
  AOI22XL U25282 ( .A0(conv_1[233]), .A1(n26059), .B0(n21623), .B1(n35231), 
        .Y(n20276) );
  OAI211XL U25283 ( .A0(n26029), .A1(n24684), .B0(n20276), .C0(n20275), .Y(
        n20280) );
  AOI22XL U25284 ( .A0(n16660), .A1(n21622), .B0(n16671), .B1(n21626), .Y(
        n20278) );
  AOI22XL U25285 ( .A0(n35195), .A1(n21627), .B0(n19179), .B1(n21624), .Y(
        n20277) );
  NAND2XL U25286 ( .A(n20278), .B(n20277), .Y(n20279) );
  AOI211XL U25287 ( .A0(n16755), .A1(n20281), .B0(n20280), .C0(n20279), .Y(
        n20282) );
  OAI211XL U25288 ( .A0(n22556), .A1(n26026), .B0(n20283), .C0(n20282), .Y(
        n20331) );
  INVXL U25289 ( .A(conv_1[236]), .Y(n31130) );
  AOI22XL U25290 ( .A0(n35195), .A1(n21687), .B0(n26081), .B1(n22599), .Y(
        n20291) );
  AOI22XL U25291 ( .A0(n19179), .A1(n21673), .B0(n16671), .B1(n21686), .Y(
        n20284) );
  OAI21XL U25292 ( .A0(n25975), .A1(n21677), .B0(n20284), .Y(n20289) );
  AOI22XL U25293 ( .A0(conv_1[221]), .A1(n26082), .B0(n34903), .B1(n22590), 
        .Y(n20286) );
  AOI22XL U25294 ( .A0(n35236), .A1(n21674), .B0(n25875), .B1(n22596), .Y(
        n20285) );
  OAI211XL U25295 ( .A0(n20287), .A1(n35159), .B0(n20286), .C0(n20285), .Y(
        n20288) );
  AOI211XL U25296 ( .A0(n16660), .A1(n21679), .B0(n20289), .C0(n20288), .Y(
        n20290) );
  OAI211XL U25297 ( .A0(n31130), .A1(n26085), .B0(n20291), .C0(n20290), .Y(
        n20330) );
  INVXL U25298 ( .A(n22490), .Y(n20292) );
  AOI221XL U25299 ( .A0(n22488), .A1(n36246), .B0(n20292), .B1(n21688), .C0(
        n28479), .Y(n20294) );
  AOI211XL U25300 ( .A0(n26081), .A1(n22487), .B0(n20294), .C0(n20293), .Y(
        n20301) );
  AOI22XL U25301 ( .A0(conv_1[220]), .A1(n26082), .B0(conv_1[235]), .B1(n26059), .Y(n20300) );
  AOI22XL U25302 ( .A0(n35195), .A1(n21644), .B0(n16671), .B1(n21651), .Y(
        n20299) );
  OAI22XL U25303 ( .A0(n21636), .A1(n18208), .B0(n21654), .B1(n35198), .Y(
        n20296) );
  OAI22XL U25304 ( .A0(n35143), .A1(n21642), .B0(n21637), .B1(n26039), .Y(
        n20295) );
  AOI211XL U25305 ( .A0(n16755), .A1(n20297), .B0(n20296), .C0(n20295), .Y(
        n20298) );
  NAND4XL U25306 ( .A(n20301), .B(n20300), .C(n20299), .D(n20298), .Y(n20329)
         );
  AOI22XL U25307 ( .A0(conv_1[234]), .A1(n26059), .B0(n26081), .B1(n22525), 
        .Y(n20310) );
  AOI22XL U25308 ( .A0(n34903), .A1(n22532), .B0(n25875), .B1(n22522), .Y(
        n20309) );
  OAI22XL U25309 ( .A0(n21659), .A1(n35239), .B0(n34543), .B1(n26029), .Y(
        n20302) );
  AOI211XL U25310 ( .A0(n26066), .A1(n22521), .B0(n20303), .C0(n20302), .Y(
        n20308) );
  OAI22XL U25311 ( .A0(n35143), .A1(n21657), .B0(n21663), .B1(n18208), .Y(
        n20305) );
  OAI22XL U25312 ( .A0(n21660), .A1(n26474), .B0(n21664), .B1(n35198), .Y(
        n20304) );
  AOI211XL U25313 ( .A0(n16755), .A1(n20306), .B0(n20305), .C0(n20304), .Y(
        n20307) );
  NAND4XL U25314 ( .A(n20310), .B(n20309), .C(n20308), .D(n20307), .Y(n20341)
         );
  NOR4XL U25315 ( .A(n20331), .B(n20330), .C(n20329), .D(n20341), .Y(n20311)
         );
  NAND4XL U25316 ( .A(n20314), .B(n20313), .C(n20312), .D(n20311), .Y(n20315)
         );
  AOI22XL U25317 ( .A0(n35236), .A1(n21757), .B0(n19179), .B1(n21755), .Y(
        n20319) );
  NAND2XL U25318 ( .A(n35195), .B(n21754), .Y(n20318) );
  OAI211XL U25319 ( .A0(n35143), .A1(n21760), .B0(n20319), .C0(n20318), .Y(
        n20326) );
  AOI22XL U25320 ( .A0(conv_1[222]), .A1(n26082), .B0(conv_1[237]), .B1(n26059), .Y(n20324) );
  AOI22XL U25321 ( .A0(n34903), .A1(n22732), .B0(n26081), .B1(n22735), .Y(
        n20323) );
  AOI22XL U25322 ( .A0(n28528), .A1(n20320), .B0(n26276), .B1(n21768), .Y(
        n20322) );
  AOI22XL U25323 ( .A0(n16660), .A1(n21775), .B0(n16671), .B1(n21767), .Y(
        n20321) );
  NAND4XL U25324 ( .A(n20324), .B(n20323), .C(n20322), .D(n20321), .Y(n20325)
         );
  AOI211XL U25325 ( .A0(n16755), .A1(n20327), .B0(n20326), .C0(n20325), .Y(
        n20328) );
  INVXL U25326 ( .A(n20328), .Y(n20343) );
  INVXL U25327 ( .A(conv_1[238]), .Y(n33846) );
  AOI22XL U25328 ( .A0(n16671), .A1(n21732), .B0(n26081), .B1(n22772), .Y(
        n20340) );
  AOI22XL U25329 ( .A0(n34903), .A1(n22771), .B0(n25879), .B1(n21735), .Y(
        n20332) );
  OAI21XL U25330 ( .A0(n20333), .A1(n26162), .B0(n20332), .Y(n20338) );
  AOI22XL U25331 ( .A0(n35195), .A1(n21727), .B0(n16660), .B1(n21728), .Y(
        n20335) );
  AOI22XL U25332 ( .A0(n35236), .A1(n21734), .B0(n19179), .B1(n21733), .Y(
        n20334) );
  OAI211XL U25333 ( .A0(n20336), .A1(n35159), .B0(n20335), .C0(n20334), .Y(
        n20337) );
  AOI211XL U25334 ( .A0(conv_1[223]), .A1(n26082), .B0(n20338), .C0(n20337), 
        .Y(n20339) );
  OAI211XL U25335 ( .A0(n33846), .A1(n26085), .B0(n20340), .C0(n20339), .Y(
        n20344) );
  NAND4XL U25336 ( .A(pool[39]), .B(n20342), .C(n20341), .D(n20344), .Y(n20346) );
  NOR3XL U25337 ( .A(pool[39]), .B(n20344), .C(n20343), .Y(n20345) );
  INVXL U25338 ( .A(n35227), .Y(n35261) );
  NAND2XL U25339 ( .A(n34844), .B(pool[35]), .Y(n20350) );
  OAI21XL U25340 ( .A0(n20351), .A1(n34844), .B0(n20350), .Y(N29251) );
  ADDFX1 U25341 ( .A(DP_OP_5170J1_126_4278_n34), .B(DP_OP_5170J1_126_4278_n38), 
        .CI(n20352), .CO(n22089), .S(n20110) );
  AOI22XL U25342 ( .A0(affine_2[27]), .A1(n33367), .B0(n16674), .B1(n20353), 
        .Y(n20354) );
  NAND2XL U25343 ( .A(n20354), .B(n33350), .Y(n16534) );
  AOI22XL U25344 ( .A0(affine_2[43]), .A1(n33367), .B0(n16674), .B1(n20356), 
        .Y(n20357) );
  NAND2XL U25345 ( .A(n20357), .B(n33340), .Y(n16550) );
  NAND2XL U25346 ( .A(counter[4]), .B(n20599), .Y(n20362) );
  INVXL U25347 ( .A(weight_2[48]), .Y(n20404) );
  OAI22XL U25348 ( .A0(n20419), .A1(n20417), .B0(n20416), .B1(n20404), .Y(
        n14644) );
  OAI22XL U25349 ( .A0(n20419), .A1(n20364), .B0(n20375), .B1(n20416), .Y(
        n14597) );
  OAI22XL U25350 ( .A0(n20419), .A1(n20366), .B0(n20365), .B1(n20416), .Y(
        n14595) );
  OAI22XL U25351 ( .A0(n20419), .A1(n20365), .B0(n20364), .B1(n20416), .Y(
        n14596) );
  OAI22XL U25352 ( .A0(n20419), .A1(n20368), .B0(n20366), .B1(n20416), .Y(
        n14594) );
  OAI22XL U25353 ( .A0(n20419), .A1(n20367), .B0(n20369), .B1(n20416), .Y(
        n14592) );
  OAI22XL U25354 ( .A0(n20419), .A1(n20369), .B0(n20368), .B1(n20416), .Y(
        n14593) );
  OAI22XL U25355 ( .A0(n20419), .A1(n20371), .B0(n20370), .B1(n20416), .Y(
        n14607) );
  INVXL U25356 ( .A(weight_2[52]), .Y(n20382) );
  OAI22XL U25357 ( .A0(n20419), .A1(n20370), .B0(n20382), .B1(n20416), .Y(
        n14608) );
  OAI22XL U25358 ( .A0(n20419), .A1(n20373), .B0(n20372), .B1(n20416), .Y(
        n14605) );
  OAI22XL U25359 ( .A0(n20419), .A1(n20372), .B0(n20371), .B1(n20416), .Y(
        n14606) );
  OAI22XL U25360 ( .A0(n20419), .A1(n20376), .B0(n20374), .B1(n20416), .Y(
        n14603) );
  OAI22XL U25361 ( .A0(n20419), .A1(n20383), .B0(n20381), .B1(n20416), .Y(
        n14611) );
  OAI22XL U25362 ( .A0(n20419), .A1(n20374), .B0(n20373), .B1(n20416), .Y(
        n14604) );
  OAI22XL U25363 ( .A0(n20419), .A1(n20375), .B0(n20377), .B1(n20416), .Y(
        n14598) );
  OAI22XL U25364 ( .A0(n20419), .A1(n20386), .B0(n20376), .B1(n20416), .Y(
        n14602) );
  INVXL U25365 ( .A(weight_2[53]), .Y(n20379) );
  OAI22XL U25366 ( .A0(n20419), .A1(n20377), .B0(n20379), .B1(n20416), .Y(
        n14599) );
  OAI22XL U25367 ( .A0(n20419), .A1(n20380), .B0(n20378), .B1(n20416), .Y(
        n14613) );
  OAI22XL U25368 ( .A0(n20419), .A1(n20378), .B0(n20385), .B1(n20416), .Y(
        n14614) );
  OAI22XL U25369 ( .A0(n20419), .A1(n20379), .B0(n36151), .B1(n20416), .Y(
        n14600) );
  OAI22XL U25370 ( .A0(n20419), .A1(n20381), .B0(n20380), .B1(n20416), .Y(
        n14612) );
  OAI22XL U25371 ( .A0(n20419), .A1(n20382), .B0(n36148), .B1(n20416), .Y(
        n14609) );
  OAI22XL U25372 ( .A0(n20419), .A1(n20384), .B0(n20383), .B1(n20416), .Y(
        n14610) );
  OAI22XL U25373 ( .A0(n20419), .A1(n20385), .B0(n20388), .B1(n20416), .Y(
        n14615) );
  OAI22XL U25374 ( .A0(n20419), .A1(n20387), .B0(n20386), .B1(n20416), .Y(
        n14601) );
  OAI22XL U25375 ( .A0(n20419), .A1(n20388), .B0(n20389), .B1(n20416), .Y(
        n14616) );
  OAI22XL U25376 ( .A0(n20419), .A1(n20396), .B0(n20399), .B1(n20416), .Y(
        n14624) );
  INVXL U25377 ( .A(weight_2[51]), .Y(n20390) );
  OAI22XL U25378 ( .A0(n20419), .A1(n20389), .B0(n20390), .B1(n20416), .Y(
        n14617) );
  OAI22XL U25379 ( .A0(n20419), .A1(n20390), .B0(n36145), .B1(n20416), .Y(
        n14618) );
  OAI22XL U25380 ( .A0(n20419), .A1(n20409), .B0(n20406), .B1(n20416), .Y(
        n14633) );
  OAI22XL U25381 ( .A0(n20419), .A1(n20391), .B0(n20392), .B1(n20416), .Y(
        n14619) );
  INVXL U25382 ( .A(weight_2[49]), .Y(n20415) );
  OAI22XL U25383 ( .A0(n20419), .A1(n20405), .B0(n20415), .B1(n20416), .Y(
        n14635) );
  OAI22XL U25384 ( .A0(n20419), .A1(n20392), .B0(n20394), .B1(n20416), .Y(
        n14620) );
  OAI22XL U25385 ( .A0(n20419), .A1(n20393), .B0(n20398), .B1(n20416), .Y(
        n14637) );
  OAI22XL U25386 ( .A0(n20419), .A1(n20394), .B0(n20395), .B1(n20416), .Y(
        n14621) );
  OAI22XL U25387 ( .A0(n20419), .A1(n20395), .B0(n20397), .B1(n20416), .Y(
        n14622) );
  OAI22XL U25388 ( .A0(n20419), .A1(n20397), .B0(n20396), .B1(n20416), .Y(
        n14623) );
  OAI22XL U25389 ( .A0(n20419), .A1(n20398), .B0(n20411), .B1(n20416), .Y(
        n14638) );
  OAI22XL U25390 ( .A0(n20419), .A1(n20399), .B0(n20400), .B1(n20416), .Y(
        n14625) );
  INVXL U25391 ( .A(weight_2[50]), .Y(n20401) );
  OAI22XL U25392 ( .A0(n20419), .A1(n20400), .B0(n20401), .B1(n20416), .Y(
        n14626) );
  OAI22XL U25393 ( .A0(n20419), .A1(n20401), .B0(n36142), .B1(n20416), .Y(
        n14627) );
  OAI22XL U25394 ( .A0(n20419), .A1(n20402), .B0(n20403), .B1(n20416), .Y(
        n14628) );
  OAI22XL U25395 ( .A0(n20419), .A1(n20403), .B0(n20407), .B1(n20416), .Y(
        n14629) );
  OAI22XL U25396 ( .A0(n20419), .A1(n20404), .B0(n36124), .B1(n20416), .Y(
        n14645) );
  OAI22XL U25397 ( .A0(n20419), .A1(n20406), .B0(n20405), .B1(n20416), .Y(
        n14634) );
  OAI22XL U25398 ( .A0(n20419), .A1(n20407), .B0(n20408), .B1(n20416), .Y(
        n14630) );
  OAI22XL U25399 ( .A0(n20419), .A1(n20408), .B0(n20410), .B1(n20416), .Y(
        n14631) );
  OAI22XL U25400 ( .A0(n20419), .A1(n20413), .B0(n20418), .B1(n20416), .Y(
        n14642) );
  OAI22XL U25401 ( .A0(n20419), .A1(n20410), .B0(n20409), .B1(n20416), .Y(
        n14632) );
  OAI22XL U25402 ( .A0(n20419), .A1(n20411), .B0(n20412), .B1(n20416), .Y(
        n14639) );
  OAI22XL U25403 ( .A0(n20419), .A1(n20412), .B0(n20414), .B1(n20416), .Y(
        n14640) );
  OAI22XL U25404 ( .A0(n20419), .A1(n20414), .B0(n20413), .B1(n20416), .Y(
        n14641) );
  OAI22XL U25405 ( .A0(n20419), .A1(n20415), .B0(n36139), .B1(n20416), .Y(
        n14636) );
  OAI22XL U25406 ( .A0(n20419), .A1(n20418), .B0(n20417), .B1(n20416), .Y(
        n14643) );
  INVXL U25407 ( .A(pool[99]), .Y(n20598) );
  AOI22XL U25408 ( .A0(n34952), .A1(n21124), .B0(n21132), .B1(n24056), .Y(
        n20421) );
  NAND2XL U25409 ( .A(n28556), .B(n21126), .Y(n20420) );
  OAI211XL U25410 ( .A0(n20422), .A1(n21959), .B0(n20421), .C0(n20420), .Y(
        n20428) );
  AOI22XL U25411 ( .A0(conv_3[228]), .A1(n21999), .B0(n22011), .B1(n21130), 
        .Y(n20426) );
  AOI2BB2XL U25412 ( .B0(conv_3[213]), .B1(n16744), .A0N(n21960), .A1N(n21123), 
        .Y(n20425) );
  AOI22XL U25413 ( .A0(n34961), .A1(n21133), .B0(n35234), .B1(n21125), .Y(
        n20424) );
  NAND4XL U25414 ( .A(n20426), .B(n20425), .C(n20424), .D(n20423), .Y(n20427)
         );
  INVXL U25415 ( .A(pool[97]), .Y(n34977) );
  AOI22XL U25416 ( .A0(conv_3[212]), .A1(n16744), .B0(n21833), .B1(n21174), 
        .Y(n20440) );
  AOI22XL U25417 ( .A0(n16667), .A1(n21169), .B0(n34961), .B1(n21176), .Y(
        n20431) );
  NAND2XL U25418 ( .A(conv_3[227]), .B(n21999), .Y(n20430) );
  OAI211XL U25419 ( .A0(n20432), .A1(n21960), .B0(n20431), .C0(n20430), .Y(
        n20438) );
  AOI22XL U25420 ( .A0(n28414), .A1(n21177), .B0(n35234), .B1(n21168), .Y(
        n20435) );
  AOI22XL U25421 ( .A0(n26376), .A1(n20433), .B0(n34954), .B1(n21170), .Y(
        n20434) );
  OAI211XL U25422 ( .A0(n20436), .A1(n35135), .B0(n20435), .C0(n20434), .Y(
        n20437) );
  AOI22XL U25423 ( .A0(n35236), .A1(n20442), .B0(n24056), .B1(n21155), .Y(
        n20444) );
  NAND2XL U25424 ( .A(n28528), .B(n21151), .Y(n20443) );
  OAI211XL U25425 ( .A0(n21148), .A1(n21960), .B0(n20444), .C0(n20443), .Y(
        n20450) );
  AOI22XL U25426 ( .A0(conv_3[211]), .A1(n16744), .B0(n22011), .B1(n21150), 
        .Y(n20448) );
  AOI22XL U25427 ( .A0(conv_3[226]), .A1(n21999), .B0(n34952), .B1(n21144), 
        .Y(n20447) );
  AOI22XL U25428 ( .A0(n34961), .A1(n21157), .B0(n35234), .B1(n21156), .Y(
        n20445) );
  NAND4XL U25429 ( .A(n20448), .B(n20447), .C(n20446), .D(n20445), .Y(n20449)
         );
  AOI222XL U25430 ( .A0(pool[95]), .A1(pool[96]), .B0(pool[95]), .B1(n34975), 
        .C0(pool[96]), .C1(n34975), .Y(n20452) );
  AOI222XL U25431 ( .A0(n34977), .A1(n34976), .B0(n34977), .B1(n20452), .C0(
        n34976), .C1(n20452), .Y(n20453) );
  AOI222XL U25432 ( .A0(n34980), .A1(pool[98]), .B0(n34980), .B1(n20453), .C0(
        pool[98]), .C1(n20453), .Y(n20537) );
  AOI22XL U25433 ( .A0(n34961), .A1(n21257), .B0(n35234), .B1(n21259), .Y(
        n20455) );
  NAND2XL U25434 ( .A(n28528), .B(n21258), .Y(n20454) );
  OAI211XL U25435 ( .A0(n19767), .A1(n21262), .B0(n20455), .C0(n20454), .Y(
        n20461) );
  AOI22XL U25436 ( .A0(n22011), .A1(n21265), .B0(n34950), .B1(n21269), .Y(
        n20459) );
  AOI22XL U25437 ( .A0(conv_3[231]), .A1(n21999), .B0(conv_3[216]), .B1(n16744), .Y(n20458) );
  AOI22XL U25438 ( .A0(n21998), .A1(n21263), .B0(n34952), .B1(n21270), .Y(
        n20457) );
  NAND4XL U25439 ( .A(n20459), .B(n20458), .C(n20457), .D(n20456), .Y(n20460)
         );
  AOI211XL U25440 ( .A0(n28465), .A1(n20462), .B0(n20461), .C0(n20460), .Y(
        n20533) );
  AOI22XL U25441 ( .A0(n35234), .A1(n21211), .B0(n34950), .B1(n21213), .Y(
        n20464) );
  NAND2XL U25442 ( .A(conv_3[232]), .B(n21999), .Y(n20463) );
  OAI211XL U25443 ( .A0(n19767), .A1(n21216), .B0(n20464), .C0(n20463), .Y(
        n20470) );
  AOI22XL U25444 ( .A0(conv_3[217]), .A1(n16744), .B0(n22011), .B1(n21228), 
        .Y(n20468) );
  AOI22XL U25445 ( .A0(n34952), .A1(n21217), .B0(n21998), .B1(n21226), .Y(
        n20467) );
  AOI22XL U25446 ( .A0(n28528), .A1(n21218), .B0(n16667), .B1(n21225), .Y(
        n20465) );
  NAND4XL U25447 ( .A(n20468), .B(n20467), .C(n20466), .D(n20465), .Y(n20469)
         );
  AOI211XL U25448 ( .A0(n28465), .A1(n20471), .B0(n20470), .C0(n20469), .Y(
        n20532) );
  NAND4XL U25449 ( .A(n20581), .B(n20588), .C(n20577), .D(n20578), .Y(n20489)
         );
  AOI22XL U25450 ( .A0(conv_3[221]), .A1(n16744), .B0(n34952), .B1(n21314), 
        .Y(n20479) );
  AOI22XL U25451 ( .A0(n16659), .A1(n21320), .B0(n24056), .B1(n21305), .Y(
        n20478) );
  OAI22XL U25452 ( .A0(n21310), .A1(n35196), .B0(n21317), .B1(n28577), .Y(
        n20475) );
  AOI22XL U25453 ( .A0(conv_3[236]), .A1(n21999), .B0(n22011), .B1(n21318), 
        .Y(n20472) );
  OAI21XL U25454 ( .A0(n20473), .A1(n21960), .B0(n20472), .Y(n20474) );
  AOI211XL U25455 ( .A0(n35236), .A1(n20476), .B0(n20475), .C0(n20474), .Y(
        n20477) );
  NAND4XL U25456 ( .A(n20480), .B(n20479), .C(n20478), .D(n20477), .Y(n20574)
         );
  AOI22XL U25457 ( .A0(n34961), .A1(n21361), .B0(n24056), .B1(n21363), .Y(
        n20488) );
  AOI22XL U25458 ( .A0(conv_3[235]), .A1(n21999), .B0(n34952), .B1(n21353), 
        .Y(n20487) );
  AOI22XL U25459 ( .A0(n35236), .A1(n20481), .B0(n22011), .B1(n21371), .Y(
        n20486) );
  OAI22XL U25460 ( .A0(n21352), .A1(n35196), .B0(n21356), .B1(n28479), .Y(
        n20484) );
  OAI21XL U25461 ( .A0(n21359), .A1(n21960), .B0(n20482), .Y(n20483) );
  AOI211XL U25462 ( .A0(n16667), .A1(n21364), .B0(n20484), .C0(n20483), .Y(
        n20485) );
  NAND4XL U25463 ( .A(n20488), .B(n20487), .C(n20486), .D(n20485), .Y(n20575)
         );
  AOI211XL U25464 ( .A0(n28465), .A1(n20489), .B0(n20574), .C0(n20575), .Y(
        n20530) );
  OAI22XL U25465 ( .A0(n20492), .A1(n20491), .B0(n23627), .B1(n22030), .Y(
        n20493) );
  AOI211XL U25466 ( .A0(n34952), .A1(n21201), .B0(n20494), .C0(n20493), .Y(
        n20502) );
  AOI22XL U25467 ( .A0(n28528), .A1(n21196), .B0(n28556), .B1(n21197), .Y(
        n20501) );
  AOI22XL U25468 ( .A0(n34961), .A1(n21190), .B0(n21202), .B1(n24056), .Y(
        n20500) );
  OAI22XL U25469 ( .A0(n20495), .A1(n21959), .B0(n22168), .B1(n22008), .Y(
        n20497) );
  OAI22XL U25470 ( .A0(n21193), .A1(n35196), .B0(n21192), .B1(n28575), .Y(
        n20496) );
  AOI211XL U25471 ( .A0(n28465), .A1(n20498), .B0(n20497), .C0(n20496), .Y(
        n20499) );
  NAND4XL U25472 ( .A(n20502), .B(n20501), .C(n20500), .D(n20499), .Y(n20531)
         );
  AOI22XL U25473 ( .A0(conv_3[230]), .A1(n21999), .B0(n22011), .B1(n21235), 
        .Y(n20512) );
  AOI22XL U25474 ( .A0(conv_3[215]), .A1(n16744), .B0(n34952), .B1(n20503), 
        .Y(n20511) );
  OAI22XL U25475 ( .A0(n21243), .A1(n18196), .B0(n21253), .B1(n35196), .Y(
        n20504) );
  OAI22XL U25476 ( .A0(n21236), .A1(n21960), .B0(n21242), .B1(n21959), .Y(
        n20507) );
  OAI22XL U25477 ( .A0(n19767), .A1(n21246), .B0(n21244), .B1(n28577), .Y(
        n20506) );
  AOI211XL U25478 ( .A0(n28465), .A1(n20508), .B0(n20507), .C0(n20506), .Y(
        n20509) );
  NAND4XL U25479 ( .A(n20512), .B(n20511), .C(n20510), .D(n20509), .Y(n20534)
         );
  AOI22XL U25480 ( .A0(n16659), .A1(n21336), .B0(n16667), .B1(n21335), .Y(
        n20520) );
  AOI22XL U25481 ( .A0(n34952), .A1(n21340), .B0(n22011), .B1(n21333), .Y(
        n20518) );
  OAI22XL U25482 ( .A0(n20513), .A1(n21959), .B0(n35675), .B1(n22008), .Y(
        n20517) );
  OAI22XL U25483 ( .A0(n20514), .A1(n21960), .B0(n32061), .B1(n22030), .Y(
        n20516) );
  OAI22XL U25484 ( .A0(n19767), .A1(n21343), .B0(n21339), .B1(n18196), .Y(
        n20515) );
  NOR4BXL U25485 ( .AN(n20518), .B(n20517), .C(n20516), .D(n20515), .Y(n20519)
         );
  NAND3XL U25486 ( .A(n20521), .B(n20520), .C(n20519), .Y(n20584) );
  AOI22XL U25487 ( .A0(n28528), .A1(n21304), .B0(n16667), .B1(n21288), .Y(
        n20528) );
  AOI22XL U25488 ( .A0(n22011), .A1(n21297), .B0(n34952), .B1(n21282), .Y(
        n20527) );
  AOI22XL U25489 ( .A0(conv_3[219]), .A1(n16744), .B0(n21998), .B1(n21295), 
        .Y(n20526) );
  OAI22XL U25490 ( .A0(n19767), .A1(n21289), .B0(n21290), .B1(n28575), .Y(
        n20524) );
  AOI22XL U25491 ( .A0(conv_3[234]), .A1(n21999), .B0(n34950), .B1(n21286), 
        .Y(n20522) );
  OAI21XL U25492 ( .A0(n21285), .A1(n35196), .B0(n20522), .Y(n20523) );
  AOI211XL U25493 ( .A0(n34961), .A1(n21287), .B0(n20524), .C0(n20523), .Y(
        n20525) );
  NAND4XL U25494 ( .A(n20528), .B(n20527), .C(n20526), .D(n20525), .Y(n20573)
         );
  NOR4XL U25495 ( .A(n20531), .B(n20534), .C(n20584), .D(n20573), .Y(n20529)
         );
  NAND4XL U25496 ( .A(n20533), .B(n20532), .C(n20530), .D(n20529), .Y(n20536)
         );
  INVXL U25497 ( .A(n20531), .Y(n20597) );
  OAI22XL U25498 ( .A0(n33904), .A1(n22008), .B0(n32142), .B1(n22030), .Y(
        n20539) );
  AOI211XL U25499 ( .A0(n22011), .A1(n20541), .B0(n20540), .C0(n20539), .Y(
        n20549) );
  AOI22XL U25500 ( .A0(n35236), .A1(n20542), .B0(n34952), .B1(n21381), .Y(
        n20548) );
  AOI22XL U25501 ( .A0(n28414), .A1(n21392), .B0(n34961), .B1(n21387), .Y(
        n20547) );
  OAI22XL U25502 ( .A0(n19767), .A1(n21385), .B0(n21393), .B1(n35196), .Y(
        n20544) );
  OAI22XL U25503 ( .A0(n21389), .A1(n28479), .B0(n21390), .B1(n28577), .Y(
        n20543) );
  AOI211XL U25504 ( .A0(n28465), .A1(n20545), .B0(n20544), .C0(n20543), .Y(
        n20546) );
  NAND4XL U25505 ( .A(n20549), .B(n20548), .C(n20547), .D(n20546), .Y(n20594)
         );
  INVXL U25506 ( .A(conv_3[223]), .Y(n32136) );
  OAI22XL U25507 ( .A0(n26274), .A1(n20550), .B0(n32136), .B1(n22030), .Y(
        n20551) );
  AOI211XL U25508 ( .A0(n22011), .A1(n21410), .B0(n20552), .C0(n20551), .Y(
        n20561) );
  AOI22XL U25509 ( .A0(n16659), .A1(n21404), .B0(n24056), .B1(n21409), .Y(
        n20560) );
  AOI22XL U25510 ( .A0(n16667), .A1(n21405), .B0(n34961), .B1(n21411), .Y(
        n20559) );
  OAI22XL U25511 ( .A0(n20554), .A1(n21960), .B0(n20553), .B1(n21959), .Y(
        n20556) );
  OAI22XL U25512 ( .A0(n21408), .A1(n28575), .B0(n21407), .B1(n35196), .Y(
        n20555) );
  AOI211XL U25513 ( .A0(n28465), .A1(n20557), .B0(n20556), .C0(n20555), .Y(
        n20558) );
  NAND4XL U25514 ( .A(n20561), .B(n20560), .C(n20559), .D(n20558), .Y(n20582)
         );
  AOI22XL U25515 ( .A0(n35236), .A1(n20562), .B0(conv_3[237]), .B1(n21999), 
        .Y(n20572) );
  AOI22XL U25516 ( .A0(n34952), .A1(n21423), .B0(n22011), .B1(n21431), .Y(
        n20571) );
  OAI22XL U25517 ( .A0(n20563), .A1(n21960), .B0(n34653), .B1(n22030), .Y(
        n20564) );
  OAI22XL U25518 ( .A0(n21433), .A1(n35196), .B0(n21428), .B1(n28479), .Y(
        n20567) );
  OAI22XL U25519 ( .A0(n21430), .A1(n28577), .B0(n21434), .B1(n18196), .Y(
        n20566) );
  AOI211XL U25520 ( .A0(n28465), .A1(n20568), .B0(n20567), .C0(n20566), .Y(
        n20569) );
  NAND4XL U25521 ( .A(n20572), .B(n20571), .C(n20570), .D(n20569), .Y(n20580)
         );
  NOR3XL U25522 ( .A(pool[99]), .B(n20582), .C(n20580), .Y(n20593) );
  INVXL U25523 ( .A(n20573), .Y(n20579) );
  INVXL U25524 ( .A(n20574), .Y(n20576) );
  INVXL U25525 ( .A(n20575), .Y(n20587) );
  NOR4BXL U25526 ( .AN(n20584), .B(n20579), .C(n20576), .D(n20587), .Y(n20591)
         );
  AOI22XL U25527 ( .A0(n20579), .A1(n20578), .B0(n20577), .B1(n20576), .Y(
        n20590) );
  INVXL U25528 ( .A(n20581), .Y(n20583) );
  OAI211XL U25529 ( .A0(n20584), .A1(n20583), .B0(pool[99]), .C0(n20582), .Y(
        n20585) );
  AOI211XL U25530 ( .A0(n20588), .A1(n20587), .B0(n20586), .C0(n20585), .Y(
        n20589) );
  OAI211XL U25531 ( .A0(n28465), .A1(n20591), .B0(n20590), .C0(n20589), .Y(
        n20592) );
  AOI22XL U25532 ( .A0(n34978), .A1(n20598), .B0(n20597), .B1(n34979), .Y(
        N29315) );
  AOI2BB1X1 U25533 ( .A0N(n20602), .A1N(n20604), .B0(n30350), .Y(n20603) );
  INVXL U25534 ( .A(filter_2[52]), .Y(n22055) );
  AOI22XL U25535 ( .A0(n20603), .A1(n36148), .B0(n22055), .B1(n22105), .Y(
        n14842) );
  INVXL U25536 ( .A(filter_2[51]), .Y(n22054) );
  AOI22XL U25537 ( .A0(n20603), .A1(n36145), .B0(n22054), .B1(n22105), .Y(
        n14841) );
  INVXL U25538 ( .A(filter_1[45]), .Y(n20606) );
  INVXL U25539 ( .A(filter_1[39]), .Y(n28233) );
  AOI22XL U25540 ( .A0(n20608), .A1(n20606), .B0(n28233), .B1(n28249), .Y(
        n14688) );
  INVXL U25541 ( .A(filter_1[51]), .Y(n20607) );
  AOI22XL U25542 ( .A0(n20608), .A1(n20607), .B0(n20606), .B1(n28249), .Y(
        n14689) );
  INVXL U25543 ( .A(filter_1[36]), .Y(n28228) );
  INVXL U25544 ( .A(filter_1[30]), .Y(n28220) );
  AOI22XL U25545 ( .A0(n20608), .A1(n28228), .B0(n28220), .B1(n28249), .Y(
        n14714) );
  INVXL U25546 ( .A(filter_1[28]), .Y(n28230) );
  INVXL U25547 ( .A(filter_1[22]), .Y(n28217) );
  AOI22XL U25548 ( .A0(n20608), .A1(n28230), .B0(n28217), .B1(n28249), .Y(
        n14676) );
  AOI22XL U25549 ( .A0(n20608), .A1(n36145), .B0(n20607), .B1(n28249), .Y(
        n14690) );
  INVXL U25550 ( .A(filter_1[46]), .Y(n28221) );
  INVXL U25551 ( .A(filter_1[40]), .Y(n24426) );
  AOI22XL U25552 ( .A0(n20608), .A1(n28221), .B0(n24426), .B1(n28249), .Y(
        n14679) );
  INVXL U25553 ( .A(filter_1[14]), .Y(n28234) );
  AOI22XL U25554 ( .A0(n20608), .A1(n28236), .B0(n28234), .B1(n28249), .Y(
        n14693) );
  AOI22XL U25555 ( .A0(n34844), .A1(n20610), .B0(n20609), .B1(n34840), .Y(
        N29255) );
  AOI22XL U25556 ( .A0(n34844), .A1(n20612), .B0(n20611), .B1(n34840), .Y(
        N29254) );
  AND2XL U25557 ( .A(n20645), .B(n20613), .Y(n20623) );
  INVXL U25558 ( .A(n20614), .Y(n20638) );
  AND2XL U25559 ( .A(n20624), .B(n20646), .Y(n20622) );
  AND2XL U25560 ( .A(n20619), .B(n20648), .Y(n20621) );
  AND2XL U25561 ( .A(n20645), .B(n20619), .Y(n20625) );
  ADDHXL U25562 ( .A(affine_1[22]), .B(n20623), .CO(DP_OP_5166J1_122_9881_n48), 
        .S(n20679) );
  AND2XL U25563 ( .A(n20645), .B(n20624), .Y(n20691) );
  AND2XL U25564 ( .A(n20624), .B(n20648), .Y(n20699) );
  ADDHXL U25565 ( .A(affine_1[21]), .B(n20625), .CO(n20620), .S(n20698) );
  AOI222XL U25566 ( .A0(n25069), .A1(affine_1[24]), .B0(n33563), .B1(n20626), 
        .C0(n29676), .C1(weight_1_bias_3[4]), .Y(n20627) );
  INVXL U25567 ( .A(n20627), .Y(n16497) );
  AND2XL U25568 ( .A(n20645), .B(n20628), .Y(n20633) );
  AND2XL U25569 ( .A(n20634), .B(n20646), .Y(n20632) );
  AND2XL U25570 ( .A(n20629), .B(n20648), .Y(n20631) );
  AND2XL U25571 ( .A(n20645), .B(n20629), .Y(n20635) );
  ADDHXL U25572 ( .A(affine_1[12]), .B(n20633), .CO(DP_OP_5167J1_123_9881_n48), 
        .S(n20670) );
  AND2XL U25573 ( .A(n20645), .B(n20634), .Y(n20683) );
  AND2XL U25574 ( .A(n20634), .B(n20648), .Y(n20687) );
  ADDHXL U25575 ( .A(affine_1[11]), .B(n20635), .CO(n20630), .S(n20686) );
  AOI222XL U25576 ( .A0(n25243), .A1(affine_1[14]), .B0(n33563), .B1(n20636), 
        .C0(n29676), .C1(weight_1_bias_2[4]), .Y(n20637) );
  INVXL U25577 ( .A(n20637), .Y(n16487) );
  AND2XL U25578 ( .A(n20645), .B(n20647), .Y(n20641) );
  AOI222XL U25579 ( .A0(n22250), .A1(affine_1[0]), .B0(n33563), .B1(n20639), 
        .C0(n29676), .C1(weight_1_bias_1[0]), .Y(n20640) );
  INVXL U25580 ( .A(n20640), .Y(n16513) );
  ADDHXL U25581 ( .A(affine_1[0]), .B(n20641), .CO(n20654), .S(n20639) );
  AND2XL U25582 ( .A(n20647), .B(n20648), .Y(n20653) );
  AND2XL U25583 ( .A(n20645), .B(n20649), .Y(n20650) );
  AOI222XL U25584 ( .A0(n22250), .A1(affine_1[1]), .B0(n33563), .B1(n20642), 
        .C0(n29676), .C1(weight_1_bias_1[1]), .Y(n20643) );
  INVXL U25585 ( .A(n20643), .Y(n16512) );
  AND2XL U25586 ( .A(n20645), .B(n20644), .Y(n20651) );
  AND2XL U25587 ( .A(n20647), .B(n20646), .Y(n20659) );
  AND2XL U25588 ( .A(n20649), .B(n20648), .Y(n20658) );
  ADDHXL U25589 ( .A(affine_1[1]), .B(n20650), .CO(n20657), .S(n20652) );
  ADDHXL U25590 ( .A(affine_1[2]), .B(n20651), .CO(DP_OP_5168J1_124_9881_n48), 
        .S(n20661) );
  ADDFX1 U25591 ( .A(n20654), .B(n20653), .CI(n20652), .CO(n20660), .S(n20642)
         );
  AOI222XL U25592 ( .A0(n22250), .A1(affine_1[2]), .B0(n33563), .B1(n20655), 
        .C0(n29676), .C1(weight_1_bias_1[2]), .Y(n20656) );
  INVXL U25593 ( .A(n20656), .Y(n16511) );
  ADDFX1 U25594 ( .A(n20662), .B(n20661), .CI(n20660), .CO(n20665), .S(n20655)
         );
  AOI222XL U25595 ( .A0(n22250), .A1(affine_1[3]), .B0(n33563), .B1(n20663), 
        .C0(n29676), .C1(weight_1_bias_1[3]), .Y(n20664) );
  INVXL U25596 ( .A(n20664), .Y(n16510) );
  ADDFX1 U25597 ( .A(DP_OP_5168J1_124_9881_n43), .B(n20666), .CI(n20665), .CO(
        n20706), .S(n20663) );
  AOI222XL U25598 ( .A0(n22250), .A1(affine_1[4]), .B0(n33563), .B1(n20667), 
        .C0(n29676), .C1(weight_1_bias_1[4]), .Y(n20668) );
  INVXL U25599 ( .A(n20668), .Y(n16509) );
  ADDFX1 U25600 ( .A(n20671), .B(n20670), .CI(n20669), .CO(n20674), .S(n20672)
         );
  AOI222XL U25601 ( .A0(n25243), .A1(affine_1[12]), .B0(n33563), .B1(n20672), 
        .C0(n29676), .C1(weight_1_bias_2[2]), .Y(n20673) );
  INVXL U25602 ( .A(n20673), .Y(n16489) );
  ADDFX1 U25603 ( .A(DP_OP_5167J1_123_9881_n43), .B(n20675), .CI(n20674), .CO(
        n20712), .S(n20676) );
  AOI222XL U25604 ( .A0(n25243), .A1(affine_1[13]), .B0(n33563), .B1(n20676), 
        .C0(n29676), .C1(weight_1_bias_2[3]), .Y(n20677) );
  INVXL U25605 ( .A(n20677), .Y(n16488) );
  ADDFX1 U25606 ( .A(n20680), .B(n20679), .CI(n20678), .CO(n20694), .S(n20681)
         );
  AOI222XL U25607 ( .A0(n25069), .A1(affine_1[22]), .B0(n33563), .B1(n20681), 
        .C0(n29676), .C1(weight_1_bias_3[2]), .Y(n20682) );
  INVXL U25608 ( .A(n20682), .Y(n16499) );
  ADDHXL U25609 ( .A(affine_1[10]), .B(n20683), .CO(n20688), .S(n20684) );
  AOI222XL U25610 ( .A0(n25243), .A1(affine_1[10]), .B0(n33563), .B1(n20684), 
        .C0(n29676), .C1(weight_1_bias_2[0]), .Y(n20685) );
  INVXL U25611 ( .A(n20685), .Y(n16491) );
  AOI222XL U25612 ( .A0(n25243), .A1(affine_1[11]), .B0(n33563), .B1(n20689), 
        .C0(n29676), .C1(weight_1_bias_2[1]), .Y(n20690) );
  INVXL U25613 ( .A(n20690), .Y(n16490) );
  ADDHXL U25614 ( .A(affine_1[20]), .B(n20691), .CO(n20700), .S(n20692) );
  AOI222XL U25615 ( .A0(n25069), .A1(affine_1[20]), .B0(n33563), .B1(n20692), 
        .C0(n29676), .C1(weight_1_bias_3[0]), .Y(n20693) );
  INVXL U25616 ( .A(n20693), .Y(n16501) );
  AOI222XL U25617 ( .A0(n25069), .A1(affine_1[23]), .B0(n33563), .B1(n20696), 
        .C0(n29676), .C1(weight_1_bias_3[3]), .Y(n20697) );
  INVXL U25618 ( .A(n20697), .Y(n16498) );
  AOI222XL U25619 ( .A0(n25069), .A1(affine_1[21]), .B0(n33563), .B1(n20701), 
        .C0(n29676), .C1(weight_1_bias_3[1]), .Y(n20702) );
  INVXL U25620 ( .A(n20702), .Y(n16500) );
  ADDFX1 U25621 ( .A(DP_OP_5166J1_122_9881_n36), .B(DP_OP_5166J1_122_9881_n42), 
        .CI(n20703), .CO(n20709), .S(n20626) );
  AOI22XL U25622 ( .A0(n33563), .A1(n20704), .B0(affine_1[26]), .B1(n25069), 
        .Y(n20705) );
  NAND2XL U25623 ( .A(n20705), .B(n33412), .Y(n16495) );
  ADDFX1 U25624 ( .A(DP_OP_5168J1_124_9881_n36), .B(DP_OP_5168J1_124_9881_n42), 
        .CI(n20706), .CO(n20715), .S(n20667) );
  AOI22XL U25625 ( .A0(n33563), .A1(n20707), .B0(affine_1[5]), .B1(n22250), 
        .Y(n20708) );
  NAND2XL U25626 ( .A(n20708), .B(n33077), .Y(n16508) );
  AOI22XL U25627 ( .A0(n33563), .A1(n20710), .B0(affine_1[25]), .B1(n25069), 
        .Y(n20711) );
  NAND2XL U25628 ( .A(n20711), .B(n33412), .Y(n16496) );
  ADDFX1 U25629 ( .A(DP_OP_5167J1_123_9881_n36), .B(DP_OP_5167J1_123_9881_n42), 
        .CI(n20712), .CO(n20723), .S(n20636) );
  AOI22XL U25630 ( .A0(n33563), .A1(n20713), .B0(affine_1[15]), .B1(n25243), 
        .Y(n20714) );
  NAND2XL U25631 ( .A(n20714), .B(n33564), .Y(n16486) );
  AOI22XL U25632 ( .A0(n33563), .A1(n20716), .B0(affine_1[6]), .B1(n22250), 
        .Y(n20717) );
  NAND2XL U25633 ( .A(n20717), .B(n33077), .Y(n16507) );
  AOI22XL U25634 ( .A0(affine_2[44]), .A1(n33367), .B0(n16674), .B1(n20719), 
        .Y(n20720) );
  NAND2XL U25635 ( .A(n20720), .B(n33340), .Y(n16549) );
  INVXL U25636 ( .A(pixel[1]), .Y(n35254) );
  AOI22XL U25637 ( .A0(n22896), .A1(n20721), .B0(n35254), .B1(n23672), .Y(
        N17495) );
  INVXL U25638 ( .A(pixel[13]), .Y(n20722) );
  INVXL U25639 ( .A(pixel[12]), .Y(n23674) );
  AOI22XL U25640 ( .A0(n22896), .A1(n20722), .B0(n23674), .B1(n23672), .Y(
        N17506) );
  INVXL U25641 ( .A(pixel[14]), .Y(n24401) );
  AOI22XL U25642 ( .A0(n22896), .A1(n24401), .B0(n20722), .B1(n23672), .Y(
        N17507) );
  ADDFX1 U25643 ( .A(DP_OP_5167J1_123_9881_n28), .B(DP_OP_5167J1_123_9881_n35), 
        .CI(n20723), .CO(n22196), .S(n20713) );
  AOI22XL U25644 ( .A0(n33563), .A1(n20724), .B0(affine_1[16]), .B1(n25243), 
        .Y(n20725) );
  NAND2XL U25645 ( .A(n20725), .B(n33564), .Y(n16485) );
  INVXL U25646 ( .A(conv_2[405]), .Y(n24211) );
  OAI2BB2XL U25647 ( .B0(n24211), .B1(n21536), .A0N(conv_2[420]), .A1N(n21765), 
        .Y(n20750) );
  INVXL U25648 ( .A(conv_2[15]), .Y(n24201) );
  INVXL U25649 ( .A(conv_2[0]), .Y(n24006) );
  OAI22XL U25650 ( .A0(n24201), .A1(n21729), .B0(n24006), .B1(n21730), .Y(
        n20749) );
  AND2XL U25651 ( .A(n22762), .B(conv_2[225]), .Y(n20727) );
  AOI22XL U25652 ( .A0(n20735), .A1(conv_2[255]), .B0(conv_2[240]), .B1(n18526), .Y(n24040) );
  AOI211XL U25653 ( .A0(conv_2[210]), .A1(n22759), .B0(n20727), .C0(n20732), 
        .Y(n34910) );
  AOI22XL U25654 ( .A0(n18810), .A1(conv_2[120]), .B0(n18658), .B1(conv_2[90]), 
        .Y(n20729) );
  NAND2XL U25655 ( .A(n20729), .B(n20728), .Y(n34907) );
  AOI22XL U25656 ( .A0(n16716), .A1(conv_2[300]), .B0(n22616), .B1(conv_2[270]), .Y(n20731) );
  NAND2XL U25657 ( .A(n20731), .B(n20730), .Y(n34911) );
  AOI22XL U25658 ( .A0(n28324), .A1(n34907), .B0(n16663), .B1(n34911), .Y(
        n20734) );
  AOI22XL U25659 ( .A0(n20735), .A1(conv_2[525]), .B0(conv_2[510]), .B1(n19253), .Y(n24043) );
  OAI21XL U25660 ( .A0(n20742), .A1(n20732), .B0(n22847), .Y(n20733) );
  OAI211XL U25661 ( .A0(n34910), .A1(n28575), .B0(n20734), .C0(n20733), .Y(
        n20748) );
  INVXL U25662 ( .A(n26285), .Y(n26260) );
  AOI22XL U25663 ( .A0(n20735), .A1(conv_2[495]), .B0(conv_2[480]), .B1(n19253), .Y(n24042) );
  AOI22XL U25664 ( .A0(conv_2[390]), .A1(n21749), .B0(n26260), .B1(n34904), 
        .Y(n20746) );
  INVXL U25665 ( .A(conv_2[465]), .Y(n22888) );
  INVXL U25666 ( .A(conv_2[450]), .Y(n34445) );
  AOI22XL U25667 ( .A0(n20735), .A1(n22888), .B0(n34445), .B1(n18526), .Y(
        n34902) );
  AOI22XL U25668 ( .A0(conv_2[435]), .A1(n21752), .B0(n21761), .B1(n34902), 
        .Y(n20745) );
  AOI22XL U25669 ( .A0(n25299), .A1(conv_2[150]), .B0(n16673), .B1(conv_2[195]), .Y(n20737) );
  NAND2XL U25670 ( .A(n20737), .B(n20736), .Y(n34913) );
  AOI22XL U25671 ( .A0(n25299), .A1(conv_2[30]), .B0(n16673), .B1(conv_2[75]), 
        .Y(n20739) );
  NAND2XL U25672 ( .A(n20739), .B(n20738), .Y(n34914) );
  AOI22XL U25673 ( .A0(n16665), .A1(n34913), .B0(n28559), .B1(n34914), .Y(
        n20744) );
  NAND2XL U25674 ( .A(n20741), .B(n20740), .Y(n34912) );
  INVXL U25675 ( .A(n21801), .Y(n34905) );
  AOI22XL U25676 ( .A0(n21756), .A1(n34912), .B0(n21736), .B1(n34905), .Y(
        n20743) );
  NAND4XL U25677 ( .A(n20746), .B(n20745), .C(n20744), .D(n20743), .Y(n20747)
         );
  NOR4XL U25678 ( .A(n20750), .B(n20749), .C(n20748), .D(n20747), .Y(n21091)
         );
  INVXL U25679 ( .A(conv_2[59]), .Y(n33108) );
  OAI22XL U25680 ( .A0(n19902), .A1(n33108), .B0(n18321), .B1(n32677), .Y(
        n20752) );
  INVXL U25681 ( .A(conv_2[44]), .Y(n27957) );
  OAI22XL U25682 ( .A0(n22740), .A1(n30247), .B0(n22717), .B1(n27957), .Y(
        n20751) );
  AOI22XL U25683 ( .A0(conv_2[419]), .A1(n21763), .B0(conv_2[239]), .B1(n21764), .Y(n20754) );
  AND2XL U25684 ( .A(n21688), .B(n25812), .Y(n21983) );
  NAND2XL U25685 ( .A(n28304), .B(n26162), .Y(n28372) );
  AOI22XL U25686 ( .A0(n21983), .A1(n28372), .B0(n25813), .B1(n21753), .Y(
        n20753) );
  OAI211XL U25687 ( .A0(n25822), .A1(n16672), .B0(n20754), .C0(n20753), .Y(
        n20771) );
  AOI22XL U25688 ( .A0(conv_2[29]), .A1(n21766), .B0(conv_2[404]), .B1(n21749), 
        .Y(n20770) );
  AOI22XL U25689 ( .A0(conv_2[449]), .A1(n21752), .B0(n21761), .B1(n25819), 
        .Y(n20769) );
  INVXL U25690 ( .A(conv_2[224]), .Y(n31126) );
  INVXL U25691 ( .A(conv_2[434]), .Y(n28897) );
  INVXL U25692 ( .A(n21765), .Y(n21567) );
  OAI22XL U25693 ( .A0(n31126), .A1(n21556), .B0(n28897), .B1(n21567), .Y(
        n20767) );
  INVXL U25694 ( .A(conv_2[14]), .Y(n27935) );
  OAI22XL U25695 ( .A0(n27935), .A1(n21730), .B0(n20755), .B1(n25815), .Y(
        n20766) );
  INVXL U25696 ( .A(conv_2[149]), .Y(n30239) );
  OAI22XL U25697 ( .A0(n19902), .A1(n30254), .B0(n18321), .B1(n30239), .Y(
        n20756) );
  INVXL U25698 ( .A(conv_2[344]), .Y(n29453) );
  INVXL U25699 ( .A(conv_2[359]), .Y(n29465) );
  INVXL U25700 ( .A(conv_2[389]), .Y(n28160) );
  OAI22XL U25701 ( .A0(n19902), .A1(n29465), .B0(n18321), .B1(n28160), .Y(
        n20758) );
  OAI22XL U25702 ( .A0(n25821), .A1(n26621), .B0(n25820), .B1(n21704), .Y(
        n20765) );
  INVXL U25703 ( .A(conv_2[329]), .Y(n33237) );
  OAI22XL U25704 ( .A0(n22550), .A1(n28890), .B0(n18750), .B1(n33237), .Y(
        n20760) );
  INVXL U25705 ( .A(conv_2[194]), .Y(n29958) );
  INVXL U25706 ( .A(conv_2[164]), .Y(n24535) );
  INVXL U25707 ( .A(conv_2[209]), .Y(n33040) );
  OAI22XL U25708 ( .A0(n22717), .A1(n24535), .B0(n22716), .B1(n33040), .Y(
        n20762) );
  OAI22XL U25709 ( .A0(n25814), .A1(n28349), .B0(n25823), .B1(n28553), .Y(
        n20764) );
  NOR4XL U25710 ( .A(n20767), .B(n20766), .C(n20765), .D(n20764), .Y(n20768)
         );
  NAND4BXL U25711 ( .AN(n20771), .B(n20770), .C(n20769), .D(n20768), .Y(n21088) );
  INVXL U25712 ( .A(n21736), .Y(n21759) );
  AOI22XL U25713 ( .A0(n21011), .A1(conv_2[109]), .B0(n22759), .B1(conv_2[94]), 
        .Y(n20772) );
  NAND2XL U25714 ( .A(n20773), .B(n20772), .Y(n25931) );
  AOI22XL U25715 ( .A0(n16662), .A1(conv_2[364]), .B0(n25299), .B1(conv_2[334]), .Y(n20774) );
  NAND2XL U25716 ( .A(n20775), .B(n20774), .Y(n25937) );
  AOI22XL U25717 ( .A0(n28366), .A1(n25931), .B0(n21756), .B1(n25937), .Y(
        n20779) );
  AOI22XL U25718 ( .A0(n22762), .A1(conv_2[49]), .B0(n22690), .B1(conv_2[34]), 
        .Y(n20776) );
  NAND2XL U25719 ( .A(n20777), .B(n20776), .Y(n25938) );
  NAND2XL U25720 ( .A(n18463), .B(n25938), .Y(n20778) );
  OAI211XL U25721 ( .A0(n25943), .A1(n21759), .B0(n20779), .C0(n20778), .Y(
        n20794) );
  INVXL U25722 ( .A(conv_2[409]), .Y(n28863) );
  INVXL U25723 ( .A(conv_2[214]), .Y(n28881) );
  OAI22XL U25724 ( .A0(n28863), .A1(n21536), .B0(n28881), .B1(n21556), .Y(
        n20793) );
  AOI22XL U25725 ( .A0(n22762), .A1(conv_2[289]), .B0(n16662), .B1(conv_2[304]), .Y(n20781) );
  NAND2XL U25726 ( .A(n20781), .B(n20780), .Y(n25932) );
  INVXL U25727 ( .A(n25932), .Y(n20784) );
  AOI22XL U25728 ( .A0(n34961), .A1(n25939), .B0(conv_2[4]), .B1(n21748), .Y(
        n20783) );
  AOI22XL U25729 ( .A0(n25940), .A1(n26260), .B0(n21464), .B1(n25930), .Y(
        n20782) );
  OAI211XL U25730 ( .A0(n20784), .A1(n28349), .B0(n20783), .C0(n20782), .Y(
        n20792) );
  AOI22XL U25731 ( .A0(n22847), .A1(n21863), .B0(conv_2[394]), .B1(n21749), 
        .Y(n20790) );
  AOI22XL U25732 ( .A0(conv_2[19]), .A1(n21766), .B0(conv_2[229]), .B1(n21764), 
        .Y(n20789) );
  AOI22XL U25733 ( .A0(conv_2[439]), .A1(n21752), .B0(n21678), .B1(n25930), 
        .Y(n20788) );
  AOI22XL U25734 ( .A0(n16662), .A1(conv_2[184]), .B0(n22759), .B1(conv_2[154]), .Y(n20785) );
  NAND2XL U25735 ( .A(n20786), .B(n20785), .Y(n25933) );
  AOI22XL U25736 ( .A0(n16665), .A1(n25933), .B0(conv_2[424]), .B1(n21765), 
        .Y(n20787) );
  NAND4XL U25737 ( .A(n20790), .B(n20789), .C(n20788), .D(n20787), .Y(n20791)
         );
  AOI22XL U25738 ( .A0(n22762), .A1(conv_2[353]), .B0(n22690), .B1(conv_2[338]), .Y(n20796) );
  NAND2XL U25739 ( .A(n20796), .B(n20795), .Y(n25972) );
  AOI2BB2XL U25740 ( .B0(n21756), .B1(n25972), .A0N(n25974), .A1N(n21759), .Y(
        n20809) );
  AOI22XL U25741 ( .A0(n22762), .A1(conv_2[173]), .B0(n22616), .B1(conv_2[158]), .Y(n20798) );
  NAND2XL U25742 ( .A(n20798), .B(n20797), .Y(n25970) );
  AOI22XL U25743 ( .A0(n22762), .A1(conv_2[53]), .B0(n22759), .B1(conv_2[38]), 
        .Y(n20800) );
  AOI22XL U25744 ( .A0(n16662), .A1(conv_2[68]), .B0(n18240), .B1(conv_2[83]), 
        .Y(n20799) );
  NAND2XL U25745 ( .A(n20800), .B(n20799), .Y(n25978) );
  AOI22XL U25746 ( .A0(n16665), .A1(n25970), .B0(n28559), .B1(n25978), .Y(
        n20808) );
  AOI22XL U25747 ( .A0(conv_2[8]), .A1(n21748), .B0(n21464), .B1(n25969), .Y(
        n20807) );
  AOI22XL U25748 ( .A0(n22762), .A1(conv_2[293]), .B0(n16662), .B1(conv_2[308]), .Y(n20801) );
  NAND2XL U25749 ( .A(n20802), .B(n20801), .Y(n25971) );
  INVXL U25750 ( .A(conv_2[413]), .Y(n30884) );
  INVXL U25751 ( .A(conv_2[428]), .Y(n28928) );
  OAI22XL U25752 ( .A0(n30884), .A1(n21536), .B0(n28928), .B1(n21567), .Y(
        n20805) );
  NAND2XL U25753 ( .A(n22847), .B(n21688), .Y(n21711) );
  OAI2BB2XL U25754 ( .B0(n20803), .B1(n21711), .A0N(n25969), .A1N(n21678), .Y(
        n20804) );
  AOI211XL U25755 ( .A0(n16663), .A1(n25971), .B0(n20805), .C0(n20804), .Y(
        n20806) );
  NAND4XL U25756 ( .A(n20809), .B(n20808), .C(n20807), .D(n20806), .Y(n20818)
         );
  AOI22XL U25757 ( .A0(conv_2[218]), .A1(n21762), .B0(n21761), .B1(n25976), 
        .Y(n20816) );
  AOI22XL U25758 ( .A0(conv_2[443]), .A1(n21752), .B0(conv_2[398]), .B1(n21749), .Y(n20815) );
  AOI22XL U25759 ( .A0(conv_2[23]), .A1(n21766), .B0(n26260), .B1(n20810), .Y(
        n20814) );
  AOI22XL U25760 ( .A0(n22762), .A1(conv_2[113]), .B0(n16662), .B1(conv_2[128]), .Y(n20812) );
  AOI22XL U25761 ( .A0(n25299), .A1(conv_2[98]), .B0(n18240), .B1(conv_2[143]), 
        .Y(n20811) );
  NAND2XL U25762 ( .A(n20812), .B(n20811), .Y(n25984) );
  AOI22XL U25763 ( .A0(n28324), .A1(n25984), .B0(conv_2[233]), .B1(n21764), 
        .Y(n20813) );
  NAND4XL U25764 ( .A(n20816), .B(n20815), .C(n20814), .D(n20813), .Y(n20817)
         );
  AOI22XL U25765 ( .A0(n22847), .A1(n25892), .B0(conv_2[440]), .B1(n21752), 
        .Y(n20839) );
  AOI22XL U25766 ( .A0(conv_2[5]), .A1(n21748), .B0(conv_2[215]), .B1(n21762), 
        .Y(n20838) );
  NAND2XL U25767 ( .A(n20820), .B(n20819), .Y(n25900) );
  AOI22XL U25768 ( .A0(n21756), .A1(n25900), .B0(n25898), .B1(n21753), .Y(
        n20837) );
  AOI22XL U25769 ( .A0(n16666), .A1(conv_2[170]), .B0(n25299), .B1(conv_2[155]), .Y(n20821) );
  NAND2XL U25770 ( .A(n20822), .B(n20821), .Y(n25901) );
  AOI22XL U25771 ( .A0(n21011), .A1(conv_2[110]), .B0(n16662), .B1(conv_2[125]), .Y(n20823) );
  NAND2XL U25772 ( .A(n20824), .B(n20823), .Y(n25902) );
  AOI22XL U25773 ( .A0(n25306), .A1(conv_2[290]), .B0(n25299), .B1(conv_2[275]), .Y(n20825) );
  NAND2XL U25774 ( .A(n20826), .B(n20825), .Y(n25893) );
  AOI22XL U25775 ( .A0(n28366), .A1(n25902), .B0(n16663), .B1(n25893), .Y(
        n20827) );
  OAI21XL U25776 ( .A0(n25896), .A1(n21759), .B0(n20827), .Y(n20835) );
  AOI22XL U25777 ( .A0(n25899), .A1(n26260), .B0(n21761), .B1(n25897), .Y(
        n20833) );
  AOI22XL U25778 ( .A0(conv_2[395]), .A1(n21749), .B0(conv_2[425]), .B1(n21765), .Y(n20832) );
  AOI22XL U25779 ( .A0(conv_2[410]), .A1(n21763), .B0(conv_2[230]), .B1(n21764), .Y(n20831) );
  AOI22XL U25780 ( .A0(n16662), .A1(conv_2[65]), .B0(n18658), .B1(conv_2[35]), 
        .Y(n20828) );
  NAND2XL U25781 ( .A(n20829), .B(n20828), .Y(n25903) );
  AOI22XL U25782 ( .A0(n28559), .A1(n25903), .B0(conv_2[20]), .B1(n21766), .Y(
        n20830) );
  NAND4XL U25783 ( .A(n20833), .B(n20832), .C(n20831), .D(n20830), .Y(n20834)
         );
  AOI211XL U25784 ( .A0(n16665), .A1(n25901), .B0(n20835), .C0(n20834), .Y(
        n20836) );
  NAND4XL U25785 ( .A(n20839), .B(n20838), .C(n20837), .D(n20836), .Y(n21030)
         );
  AOI22XL U25786 ( .A0(conv_2[235]), .A1(n21764), .B0(n21751), .B1(n21914), 
        .Y(n20862) );
  AOI22XL U25787 ( .A0(conv_2[445]), .A1(n21752), .B0(conv_2[430]), .B1(n21765), .Y(n20861) );
  AOI22XL U25788 ( .A0(n22616), .A1(conv_2[100]), .B0(n18240), .B1(conv_2[145]), .Y(n20841) );
  AOI22XL U25789 ( .A0(n16666), .A1(conv_2[115]), .B0(n16662), .B1(conv_2[130]), .Y(n20840) );
  NAND2XL U25790 ( .A(n20841), .B(n20840), .Y(n26036) );
  INVXL U25791 ( .A(conv_2[415]), .Y(n36040) );
  INVXL U25792 ( .A(conv_2[400]), .Y(n33140) );
  OAI22XL U25793 ( .A0(n26038), .A1(n21237), .B0(n33140), .B1(n21731), .Y(
        n20842) );
  AOI211XL U25794 ( .A0(n28324), .A1(n26036), .B0(n20843), .C0(n20842), .Y(
        n20860) );
  NAND2XL U25795 ( .A(n22713), .B(n21913), .Y(n26028) );
  NAND2XL U25796 ( .A(n26028), .B(n26037), .Y(n26033) );
  INVXL U25797 ( .A(conv_2[70]), .Y(n30124) );
  INVXL U25798 ( .A(conv_2[40]), .Y(n33590) );
  INVXL U25799 ( .A(conv_2[85]), .Y(n33816) );
  OAI22XL U25800 ( .A0(n22717), .A1(n33590), .B0(n18321), .B1(n33816), .Y(
        n20844) );
  AOI211XL U25801 ( .A0(conv_2[55]), .A1(n22762), .B0(n20845), .C0(n20844), 
        .Y(n26041) );
  AOI22XL U25802 ( .A0(n16662), .A1(conv_2[190]), .B0(n25299), .B1(conv_2[160]), .Y(n20847) );
  NAND2XL U25803 ( .A(n20847), .B(n20846), .Y(n26034) );
  AOI22XL U25804 ( .A0(n22770), .A1(conv_2[295]), .B0(n16662), .B1(conv_2[310]), .Y(n20848) );
  NAND2XL U25805 ( .A(n20849), .B(n20848), .Y(n26035) );
  AOI22XL U25806 ( .A0(n16665), .A1(n26034), .B0(n16663), .B1(n26035), .Y(
        n20852) );
  OAI2BB1XL U25807 ( .A0N(n36246), .A1N(n26032), .B0(n26028), .Y(n20850) );
  NAND2XL U25808 ( .A(n22847), .B(n20850), .Y(n20851) );
  OAI211XL U25809 ( .A0(n26041), .A1(n16672), .B0(n20852), .C0(n20851), .Y(
        n20858) );
  INVXL U25810 ( .A(conv_2[355]), .Y(n29485) );
  INVXL U25811 ( .A(conv_2[340]), .Y(n29615) );
  OAI2BB2XL U25812 ( .B0(n22717), .B1(n29615), .A0N(n16673), .A1N(conv_2[385]), 
        .Y(n20853) );
  AOI22XL U25813 ( .A0(conv_2[220]), .A1(n21762), .B0(n21678), .B1(n26032), 
        .Y(n20856) );
  AOI22XL U25814 ( .A0(conv_2[25]), .A1(n21766), .B0(conv_2[10]), .B1(n21748), 
        .Y(n20855) );
  OAI211XL U25815 ( .A0(n26040), .A1(n21704), .B0(n20856), .C0(n20855), .Y(
        n20857) );
  AOI211XL U25816 ( .A0(n21736), .A1(n26033), .B0(n20858), .C0(n20857), .Y(
        n20859) );
  NAND4XL U25817 ( .A(n20862), .B(n20861), .C(n20860), .D(n20859), .Y(n21081)
         );
  INVXL U25818 ( .A(conv_2[144]), .Y(n30093) );
  OAI22XL U25819 ( .A0(n22546), .A1(n30136), .B0(n18321), .B1(n30093), .Y(
        n20863) );
  AOI22XL U25820 ( .A0(n16662), .A1(conv_2[69]), .B0(n25299), .B1(conv_2[39]), 
        .Y(n20866) );
  AOI22XL U25821 ( .A0(n22770), .A1(conv_2[54]), .B0(n16673), .B1(conv_2[84]), 
        .Y(n20865) );
  NAND2XL U25822 ( .A(n20866), .B(n20865), .Y(n25996) );
  AOI22XL U25823 ( .A0(n22762), .A1(conv_2[294]), .B0(n22690), .B1(conv_2[279]), .Y(n20868) );
  AOI22XL U25824 ( .A0(n16662), .A1(conv_2[309]), .B0(n16673), .B1(conv_2[324]), .Y(n20867) );
  NAND2XL U25825 ( .A(n20868), .B(n20867), .Y(n25995) );
  AOI22XL U25826 ( .A0(n28559), .A1(n25996), .B0(n16663), .B1(n25995), .Y(
        n20872) );
  AOI22XL U25827 ( .A0(n16662), .A1(conv_2[369]), .B0(n22690), .B1(conv_2[339]), .Y(n20870) );
  NAND2XL U25828 ( .A(n20870), .B(n20869), .Y(n25994) );
  NAND2XL U25829 ( .A(n21756), .B(n25994), .Y(n20871) );
  OAI211XL U25830 ( .A0(n25998), .A1(n26621), .B0(n20872), .C0(n20871), .Y(
        n20886) );
  INVXL U25831 ( .A(n21751), .Y(n21712) );
  OAI22XL U25832 ( .A0(n25988), .A1(n21712), .B0(n34640), .B1(n21731), .Y(
        n20885) );
  INVXL U25833 ( .A(conv_2[159]), .Y(n34627) );
  OAI22XL U25834 ( .A0(n22612), .A1(n29893), .B0(n22717), .B1(n34627), .Y(
        n20873) );
  AOI22XL U25835 ( .A0(conv_2[444]), .A1(n21752), .B0(n21761), .B1(n25992), 
        .Y(n20877) );
  OR2XL U25836 ( .A(n36246), .B(n25997), .Y(n20875) );
  OAI2BB1XL U25837 ( .A0N(n25989), .A1N(n20875), .B0(n22847), .Y(n20876) );
  OAI211XL U25838 ( .A0(n25999), .A1(n28553), .B0(n20877), .C0(n20876), .Y(
        n20884) );
  AOI22XL U25839 ( .A0(conv_2[429]), .A1(n21765), .B0(n21678), .B1(n20878), 
        .Y(n20882) );
  AOI22XL U25840 ( .A0(conv_2[24]), .A1(n21766), .B0(conv_2[219]), .B1(n21762), 
        .Y(n20881) );
  AOI22XL U25841 ( .A0(conv_2[414]), .A1(n21763), .B0(conv_2[9]), .B1(n21748), 
        .Y(n20880) );
  AOI22XL U25842 ( .A0(conv_2[234]), .A1(n21764), .B0(n21736), .B1(n25993), 
        .Y(n20879) );
  NAND4XL U25843 ( .A(n20882), .B(n20881), .C(n20880), .D(n20879), .Y(n20883)
         );
  NOR4XL U25844 ( .A(n20886), .B(n20885), .C(n20884), .D(n20883), .Y(n21036)
         );
  AOI22XL U25845 ( .A0(n16666), .A1(conv_2[56]), .B0(n22690), .B1(conv_2[41]), 
        .Y(n20887) );
  NAND2XL U25846 ( .A(n20888), .B(n20887), .Y(n26018) );
  AOI22XL U25847 ( .A0(n28559), .A1(n26018), .B0(n21678), .B1(n26007), .Y(
        n20908) );
  OAI22XL U25848 ( .A0(n26009), .A1(n21712), .B0(n27696), .B1(n21730), .Y(
        n20907) );
  INVXL U25849 ( .A(n21711), .Y(n21725) );
  AOI22XL U25850 ( .A0(conv_2[416]), .A1(n21763), .B0(n21725), .B1(n21925), 
        .Y(n20892) );
  AOI22XL U25851 ( .A0(conv_2[26]), .A1(n21766), .B0(conv_2[401]), .B1(n21749), 
        .Y(n20891) );
  AOI22XL U25852 ( .A0(conv_2[431]), .A1(n21765), .B0(n21464), .B1(n26007), 
        .Y(n20890) );
  NAND2XL U25853 ( .A(n26015), .B(n21736), .Y(n20889) );
  NAND4XL U25854 ( .A(n20892), .B(n20891), .C(n20890), .D(n20889), .Y(n20906)
         );
  AOI22XL U25855 ( .A0(conv_2[236]), .A1(n21764), .B0(n21761), .B1(n26011), 
        .Y(n20904) );
  AOI22XL U25856 ( .A0(conv_2[446]), .A1(n21752), .B0(conv_2[221]), .B1(n21762), .Y(n20903) );
  AOI22XL U25857 ( .A0(n20978), .A1(conv_2[296]), .B0(n22616), .B1(conv_2[281]), .Y(n20893) );
  NAND2XL U25858 ( .A(n20894), .B(n20893), .Y(n26017) );
  INVXL U25859 ( .A(conv_2[146]), .Y(n34362) );
  INVXL U25860 ( .A(conv_2[116]), .Y(n34647) );
  INVXL U25861 ( .A(conv_2[101]), .Y(n30218) );
  OAI22XL U25862 ( .A0(n22546), .A1(n34647), .B0(n22717), .B1(n30218), .Y(
        n20895) );
  AOI2BB2XL U25863 ( .B0(n16663), .B1(n26017), .A0N(n26014), .A1N(n26621), .Y(
        n20902) );
  AOI22XL U25864 ( .A0(n16662), .A1(conv_2[191]), .B0(n22690), .B1(conv_2[161]), .Y(n20898) );
  NAND2XL U25865 ( .A(n20898), .B(n20897), .Y(n26008) );
  AOI22XL U25866 ( .A0(n16662), .A1(conv_2[371]), .B0(n22759), .B1(conv_2[341]), .Y(n20899) );
  NAND2XL U25867 ( .A(n20900), .B(n20899), .Y(n26016) );
  AOI22XL U25868 ( .A0(n16665), .A1(n26008), .B0(n21756), .B1(n26016), .Y(
        n20901) );
  NAND4XL U25869 ( .A(n20904), .B(n20903), .C(n20902), .D(n20901), .Y(n20905)
         );
  NOR4BXL U25870 ( .AN(n20908), .B(n20907), .C(n20906), .D(n20905), .Y(n21034)
         );
  OAI2BB1XL U25871 ( .A0N(n21004), .A1N(n21311), .B0(n25949), .Y(n20930) );
  INVXL U25872 ( .A(conv_2[426]), .Y(n28934) );
  OAI22XL U25873 ( .A0(n29086), .A1(n21729), .B0(n28934), .B1(n21567), .Y(
        n20929) );
  INVXL U25874 ( .A(conv_2[81]), .Y(n35871) );
  OAI22XL U25875 ( .A0(n22717), .A1(n27733), .B0(n18321), .B1(n35871), .Y(
        n20910) );
  INVXL U25876 ( .A(conv_2[51]), .Y(n27824) );
  OAI22XL U25877 ( .A0(n19902), .A1(n27824), .B0(n22612), .B1(n30105), .Y(
        n20909) );
  AOI22XL U25878 ( .A0(n22762), .A1(conv_2[111]), .B0(n16662), .B1(conv_2[126]), .Y(n20912) );
  NAND2XL U25879 ( .A(n20912), .B(n20911), .Y(n25952) );
  AOI22XL U25880 ( .A0(n28366), .A1(n25952), .B0(n25956), .B1(n21736), .Y(
        n20916) );
  AOI22XL U25881 ( .A0(n16662), .A1(conv_2[366]), .B0(n25299), .B1(conv_2[336]), .Y(n20914) );
  NAND2XL U25882 ( .A(n20914), .B(n20913), .Y(n25957) );
  NAND2XL U25883 ( .A(n21756), .B(n25957), .Y(n20915) );
  OAI211XL U25884 ( .A0(n25963), .A1(n16672), .B0(n20916), .C0(n20915), .Y(
        n20928) );
  INVXL U25885 ( .A(n25955), .Y(n21894) );
  AOI22XL U25886 ( .A0(conv_2[441]), .A1(n21752), .B0(n21725), .B1(n21894), 
        .Y(n20926) );
  AOI22XL U25887 ( .A0(n22762), .A1(conv_2[291]), .B0(n25299), .B1(conv_2[276]), .Y(n20917) );
  NAND2XL U25888 ( .A(n20918), .B(n20917), .Y(n25950) );
  AOI22XL U25889 ( .A0(conv_2[231]), .A1(n21764), .B0(n16663), .B1(n25950), 
        .Y(n20925) );
  AOI22XL U25890 ( .A0(conv_2[216]), .A1(n21762), .B0(n21761), .B1(n25960), 
        .Y(n20924) );
  AOI22XL U25891 ( .A0(n16662), .A1(conv_2[186]), .B0(n18240), .B1(conv_2[201]), .Y(n20920) );
  AOI22XL U25892 ( .A0(n22762), .A1(conv_2[171]), .B0(n22759), .B1(conv_2[156]), .Y(n20919) );
  NAND2XL U25893 ( .A(n20920), .B(n20919), .Y(n25951) );
  INVXL U25894 ( .A(conv_2[411]), .Y(n29491) );
  OAI22XL U25895 ( .A0(n25958), .A1(n21712), .B0(n29491), .B1(n21536), .Y(
        n20922) );
  INVXL U25896 ( .A(conv_2[396]), .Y(n28113) );
  OAI22XL U25897 ( .A0(n28113), .A1(n21731), .B0(n28777), .B1(n21730), .Y(
        n20921) );
  AOI211XL U25898 ( .A0(n16665), .A1(n25951), .B0(n20922), .C0(n20921), .Y(
        n20923) );
  NAND4XL U25899 ( .A(n20926), .B(n20925), .C(n20924), .D(n20923), .Y(n20927)
         );
  NOR4BXL U25900 ( .AN(n20930), .B(n20929), .C(n20928), .D(n20927), .Y(n21029)
         );
  AOI22XL U25901 ( .A0(n22762), .A1(conv_2[172]), .B0(n16662), .B1(conv_2[187]), .Y(n20931) );
  NAND2XL U25902 ( .A(n20932), .B(n20931), .Y(n25916) );
  AOI22XL U25903 ( .A0(n22762), .A1(conv_2[52]), .B0(n22759), .B1(conv_2[37]), 
        .Y(n20934) );
  AOI22XL U25904 ( .A0(n16662), .A1(conv_2[67]), .B0(n16673), .B1(conv_2[82]), 
        .Y(n20933) );
  NAND2XL U25905 ( .A(n20934), .B(n20933), .Y(n25920) );
  AOI22XL U25906 ( .A0(n16665), .A1(n25916), .B0(n28559), .B1(n25920), .Y(
        n20945) );
  AOI22XL U25907 ( .A0(n25299), .A1(conv_2[97]), .B0(n18240), .B1(conv_2[142]), 
        .Y(n20936) );
  AOI22XL U25908 ( .A0(n16666), .A1(conv_2[112]), .B0(n16662), .B1(conv_2[127]), .Y(n20935) );
  NAND2XL U25909 ( .A(n20936), .B(n20935), .Y(n25919) );
  AOI22XL U25910 ( .A0(n22762), .A1(conv_2[292]), .B0(n16662), .B1(conv_2[307]), .Y(n20938) );
  NAND2XL U25911 ( .A(n20938), .B(n20937), .Y(n25921) );
  AOI22XL U25912 ( .A0(n28366), .A1(n25919), .B0(n16663), .B1(n25921), .Y(
        n20944) );
  AOI22XL U25913 ( .A0(n21749), .A1(conv_2[397]), .B0(n21464), .B1(n25911), 
        .Y(n20943) );
  OAI22XL U25914 ( .A0(n20939), .A1(n21004), .B0(n25915), .B1(n21711), .Y(
        n20941) );
  INVXL U25915 ( .A(conv_2[427]), .Y(n28910) );
  INVXL U25916 ( .A(conv_2[232]), .Y(n32879) );
  OAI22XL U25917 ( .A0(n28910), .A1(n21567), .B0(n32879), .B1(n21710), .Y(
        n20940) );
  AOI211XL U25918 ( .A0(n21736), .A1(n25917), .B0(n20941), .C0(n20940), .Y(
        n20942) );
  NAND4XL U25919 ( .A(n20945), .B(n20944), .C(n20943), .D(n20942), .Y(n20954)
         );
  INVXL U25920 ( .A(n20946), .Y(n25912) );
  AOI22XL U25921 ( .A0(n21761), .A1(n25918), .B0(n21751), .B1(n25912), .Y(
        n20952) );
  AOI22XL U25922 ( .A0(conv_2[442]), .A1(n21752), .B0(conv_2[7]), .B1(n21748), 
        .Y(n20951) );
  AOI22XL U25923 ( .A0(conv_2[22]), .A1(n21766), .B0(conv_2[217]), .B1(n21762), 
        .Y(n20950) );
  AOI22XL U25924 ( .A0(n16662), .A1(conv_2[367]), .B0(n22759), .B1(conv_2[337]), .Y(n20948) );
  NAND2XL U25925 ( .A(n20948), .B(n20947), .Y(n25922) );
  AOI22XL U25926 ( .A0(conv_2[412]), .A1(n21763), .B0(n21756), .B1(n25922), 
        .Y(n20949) );
  NAND4XL U25927 ( .A(n20952), .B(n20951), .C(n20950), .D(n20949), .Y(n20953)
         );
  NAND4XL U25928 ( .A(n21036), .B(n21034), .C(n21029), .D(n21028), .Y(n20955)
         );
  NOR3XL U25929 ( .A(n21030), .B(n21081), .C(n20955), .Y(n20956) );
  AOI31XL U25930 ( .A0(n22053), .A1(n21035), .A2(n20956), .B0(pool[69]), .Y(
        n21033) );
  AOI22XL U25931 ( .A0(n16666), .A1(conv_2[48]), .B0(n16662), .B1(conv_2[63]), 
        .Y(n20957) );
  NAND2XL U25932 ( .A(n20958), .B(n20957), .Y(n25842) );
  NAND2XL U25933 ( .A(n21818), .B(n21358), .Y(n25833) );
  NAND2XL U25934 ( .A(n25833), .B(n25831), .Y(n21817) );
  AOI22XL U25935 ( .A0(n16662), .A1(conv_2[303]), .B0(n22759), .B1(conv_2[273]), .Y(n20959) );
  NAND2XL U25936 ( .A(n20960), .B(n20959), .Y(n25841) );
  AOI22XL U25937 ( .A0(n16663), .A1(n25841), .B0(n25838), .B1(n21753), .Y(
        n20961) );
  OAI21XL U25938 ( .A0(n21817), .A1(n21759), .B0(n20961), .Y(n20977) );
  AOI2BB2XL U25939 ( .B0(conv_2[18]), .B1(n21766), .A0N(n21712), .A1N(n25836), 
        .Y(n20975) );
  AOI22XL U25940 ( .A0(conv_2[408]), .A1(n21763), .B0(conv_2[3]), .B1(n21748), 
        .Y(n20974) );
  NAND2XL U25941 ( .A(n20963), .B(n20962), .Y(n25840) );
  NAND2XL U25942 ( .A(n20965), .B(n20964), .Y(n25834) );
  AOI22XL U25943 ( .A0(n16665), .A1(n25840), .B0(n28324), .B1(n25834), .Y(
        n20973) );
  AOI22XL U25944 ( .A0(n25289), .A1(conv_2[363]), .B0(n22759), .B1(conv_2[333]), .Y(n20967) );
  NAND2XL U25945 ( .A(n20967), .B(n20966), .Y(n25839) );
  AOI22XL U25946 ( .A0(conv_2[213]), .A1(n21762), .B0(n21756), .B1(n25839), 
        .Y(n20971) );
  INVXL U25947 ( .A(conv_2[393]), .Y(n29570) );
  OAI22XL U25948 ( .A0(n29558), .A1(n17171), .B0(n29570), .B1(n21731), .Y(
        n20970) );
  INVXL U25949 ( .A(conv_2[228]), .Y(n22965) );
  OAI22XL U25950 ( .A0(n22965), .A1(n21710), .B0(n32874), .B1(n21567), .Y(
        n20969) );
  OAI22XL U25951 ( .A0(n21819), .A1(n21237), .B0(n21818), .B1(n21711), .Y(
        n20968) );
  NOR4BXL U25952 ( .AN(n20971), .B(n20970), .C(n20969), .D(n20968), .Y(n20972)
         );
  NAND4XL U25953 ( .A(n20975), .B(n20974), .C(n20973), .D(n20972), .Y(n20976)
         );
  AOI22XL U25954 ( .A0(conv_2[407]), .A1(n21763), .B0(conv_2[227]), .B1(n21764), .Y(n21001) );
  AOI22XL U25955 ( .A0(conv_2[17]), .A1(n21766), .B0(conv_2[212]), .B1(n21762), 
        .Y(n21000) );
  AOI22XL U25956 ( .A0(n20978), .A1(conv_2[167]), .B0(n16662), .B1(conv_2[182]), .Y(n20979) );
  NAND2XL U25957 ( .A(n20980), .B(n20979), .Y(n25859) );
  OAI2BB1XL U25958 ( .A0N(n21688), .A1N(n20981), .B0(n20983), .Y(n25857) );
  AOI22XL U25959 ( .A0(n16665), .A1(n25859), .B0(n21736), .B1(n25857), .Y(
        n20999) );
  AOI22XL U25960 ( .A0(n21748), .A1(conv_2[2]), .B0(n21725), .B1(n20981), .Y(
        n20982) );
  OAI21XL U25961 ( .A0(n26285), .A1(n20983), .B0(n20982), .Y(n20997) );
  AOI22XL U25962 ( .A0(conv_2[437]), .A1(n21752), .B0(conv_2[392]), .B1(n21749), .Y(n20995) );
  AOI22XL U25963 ( .A0(n16662), .A1(conv_2[362]), .B0(n18658), .B1(conv_2[332]), .Y(n20985) );
  NAND2XL U25964 ( .A(n20985), .B(n20984), .Y(n25856) );
  AOI22XL U25965 ( .A0(conv_2[422]), .A1(n21765), .B0(n21756), .B1(n25856), 
        .Y(n20994) );
  NAND2XL U25966 ( .A(n20987), .B(n20986), .Y(n25860) );
  AOI22XL U25967 ( .A0(n16666), .A1(conv_2[47]), .B0(n22759), .B1(conv_2[32]), 
        .Y(n20988) );
  NAND2XL U25968 ( .A(n20989), .B(n20988), .Y(n25858) );
  AOI22XL U25969 ( .A0(n28366), .A1(n25860), .B0(n28559), .B1(n25858), .Y(
        n20993) );
  AOI22XL U25970 ( .A0(n16662), .A1(conv_2[302]), .B0(n22759), .B1(conv_2[272]), .Y(n20990) );
  NAND2XL U25971 ( .A(n20991), .B(n20990), .Y(n25850) );
  AOI22XL U25972 ( .A0(n16663), .A1(n25850), .B0(n25867), .B1(n21753), .Y(
        n20992) );
  NAND4XL U25973 ( .A(n20995), .B(n20994), .C(n20993), .D(n20992), .Y(n20996)
         );
  AOI211XL U25974 ( .A0(n21761), .A1(n25855), .B0(n20997), .C0(n20996), .Y(
        n20998) );
  NAND4XL U25975 ( .A(n21001), .B(n21000), .C(n20999), .D(n20998), .Y(n34889)
         );
  AOI22XL U25976 ( .A0(n22762), .A1(conv_2[106]), .B0(n22690), .B1(conv_2[91]), 
        .Y(n21002) );
  AOI22XL U25977 ( .A0(n28366), .A1(n25880), .B0(conv_2[16]), .B1(n21766), .Y(
        n21025) );
  NAND2XL U25978 ( .A(n22713), .B(n25874), .Y(n21848) );
  OAI22XL U25979 ( .A0(n25873), .A1(n21004), .B0(n28277), .B1(n21848), .Y(
        n21024) );
  AOI22XL U25980 ( .A0(n21761), .A1(n25876), .B0(n21751), .B1(n21849), .Y(
        n21010) );
  AOI22XL U25981 ( .A0(conv_2[406]), .A1(n21763), .B0(conv_2[226]), .B1(n21764), .Y(n21009) );
  AOI22XL U25982 ( .A0(conv_2[421]), .A1(n21765), .B0(conv_2[1]), .B1(n21748), 
        .Y(n21008) );
  AOI22XL U25983 ( .A0(n21011), .A1(conv_2[286]), .B0(n16662), .B1(conv_2[301]), .Y(n21005) );
  NAND2XL U25984 ( .A(n21006), .B(n21005), .Y(n25881) );
  NAND2XL U25985 ( .A(n16663), .B(n25881), .Y(n21007) );
  NAND4XL U25986 ( .A(n21010), .B(n21009), .C(n21008), .D(n21007), .Y(n21023)
         );
  AOI22XL U25987 ( .A0(conv_2[436]), .A1(n21752), .B0(conv_2[211]), .B1(n21762), .Y(n21021) );
  INVXL U25988 ( .A(n25873), .Y(n21845) );
  AOI22XL U25989 ( .A0(conv_2[391]), .A1(n21749), .B0(n21464), .B1(n21845), 
        .Y(n21020) );
  OAI2BB1XL U25990 ( .A0N(n36246), .A1N(n21849), .B0(n21848), .Y(n25878) );
  AOI22XL U25991 ( .A0(n16662), .A1(conv_2[361]), .B0(n22690), .B1(conv_2[331]), .Y(n21012) );
  AOI22XL U25992 ( .A0(n21736), .A1(n25878), .B0(n21756), .B1(n25882), .Y(
        n21019) );
  AOI22XL U25993 ( .A0(n16662), .A1(conv_2[181]), .B0(n16673), .B1(conv_2[196]), .Y(n21015) );
  AOI22XL U25994 ( .A0(n22762), .A1(conv_2[46]), .B0(n22690), .B1(conv_2[31]), 
        .Y(n21017) );
  NAND2XL U25995 ( .A(n21017), .B(n21016), .Y(n25877) );
  AOI22XL U25996 ( .A0(n16665), .A1(n25870), .B0(n18463), .B1(n25877), .Y(
        n21018) );
  NAND4XL U25997 ( .A(n21021), .B(n21020), .C(n21019), .D(n21018), .Y(n21022)
         );
  AOI222XL U25998 ( .A0(pool[65]), .A1(pool[66]), .B0(pool[65]), .B1(n34887), 
        .C0(pool[66]), .C1(n34887), .Y(n21026) );
  AOI222XL U25999 ( .A0(n34891), .A1(n34889), .B0(n34891), .B1(n21026), .C0(
        n34889), .C1(n21026), .Y(n21027) );
  AOI222XL U26000 ( .A0(n22051), .A1(pool[68]), .B0(n22051), .B1(n21027), .C0(
        pool[68]), .C1(n21027), .Y(n21032) );
  NOR4XL U26001 ( .A(n21036), .B(n21035), .C(n21034), .D(n22052), .Y(n21082)
         );
  AOI22XL U26002 ( .A0(conv_2[222]), .A1(n21762), .B0(n21761), .B1(n26067), 
        .Y(n21058) );
  NAND2XL U26003 ( .A(n22765), .B(n21997), .Y(n26063) );
  AOI2BB2XL U26004 ( .B0(conv_2[447]), .B1(n21752), .A0N(n28277), .A1N(n26063), 
        .Y(n21057) );
  AOI22XL U26005 ( .A0(n16716), .A1(conv_2[312]), .B0(n16673), .B1(conv_2[327]), .Y(n21038) );
  AOI22XL U26006 ( .A0(n22347), .A1(conv_2[297]), .B0(n22759), .B1(conv_2[282]), .Y(n21037) );
  NAND2XL U26007 ( .A(n21038), .B(n21037), .Y(n26058) );
  NAND2XL U26008 ( .A(n21040), .B(n21039), .Y(n26060) );
  AOI22XL U26009 ( .A0(n16663), .A1(n26058), .B0(n21756), .B1(n26060), .Y(
        n21056) );
  AOI22XL U26010 ( .A0(conv_2[237]), .A1(n21764), .B0(conv_2[417]), .B1(n21763), .Y(n21041) );
  OAI21XL U26011 ( .A0(n26285), .A1(n21046), .B0(n21041), .Y(n21054) );
  AOI22XL U26012 ( .A0(conv_2[27]), .A1(n21766), .B0(conv_2[402]), .B1(n21749), 
        .Y(n21052) );
  NAND2XL U26013 ( .A(n21043), .B(n21042), .Y(n26069) );
  AOI22XL U26014 ( .A0(n28559), .A1(n26069), .B0(conv_2[432]), .B1(n21765), 
        .Y(n21051) );
  NAND2XL U26015 ( .A(n21045), .B(n21044), .Y(n26071) );
  NAND2XL U26016 ( .A(n26063), .B(n21046), .Y(n26070) );
  AOI22XL U26017 ( .A0(n16665), .A1(n26071), .B0(n21736), .B1(n26070), .Y(
        n21050) );
  AOI22XL U26018 ( .A0(n16662), .A1(conv_2[132]), .B0(n22759), .B1(conv_2[102]), .Y(n21048) );
  AOI22XL U26019 ( .A0(n22347), .A1(conv_2[117]), .B0(n16673), .B1(conv_2[147]), .Y(n21047) );
  NAND2XL U26020 ( .A(n21048), .B(n21047), .Y(n26068) );
  AOI22XL U26021 ( .A0(n28324), .A1(n26068), .B0(n26064), .B1(n21753), .Y(
        n21049) );
  NAND4XL U26022 ( .A(n21052), .B(n21051), .C(n21050), .D(n21049), .Y(n21053)
         );
  AOI211XL U26023 ( .A0(conv_2[12]), .A1(n21748), .B0(n21054), .C0(n21053), 
        .Y(n21055) );
  NAND4XL U26024 ( .A(n21058), .B(n21057), .C(n21056), .D(n21055), .Y(n21084)
         );
  NAND2XL U26025 ( .A(n22743), .B(n21059), .Y(n26083) );
  AOI22XL U26026 ( .A0(n22847), .A1(n22027), .B0(conv_2[448]), .B1(n21752), 
        .Y(n21080) );
  AOI22XL U26027 ( .A0(conv_2[28]), .A1(n21766), .B0(conv_2[13]), .B1(n21748), 
        .Y(n21079) );
  AOI22XL U26028 ( .A0(n22347), .A1(conv_2[178]), .B0(n25299), .B1(conv_2[163]), .Y(n21061) );
  AOI22XL U26029 ( .A0(n16662), .A1(conv_2[193]), .B0(n18240), .B1(conv_2[208]), .Y(n21060) );
  NAND2XL U26030 ( .A(n21061), .B(n21060), .Y(n26091) );
  AOI22XL U26031 ( .A0(n16662), .A1(conv_2[373]), .B0(n18658), .B1(conv_2[343]), .Y(n21063) );
  NAND2XL U26032 ( .A(n21063), .B(n21062), .Y(n26092) );
  AOI22XL U26033 ( .A0(n16665), .A1(n26091), .B0(n21756), .B1(n26092), .Y(
        n21078) );
  NAND2XL U26034 ( .A(n21065), .B(n21064), .Y(n26093) );
  INVXL U26035 ( .A(conv_2[148]), .Y(n30233) );
  INVXL U26036 ( .A(conv_2[118]), .Y(n30248) );
  INVXL U26037 ( .A(conv_2[103]), .Y(n33292) );
  OAI22XL U26038 ( .A0(n19902), .A1(n30248), .B0(n22717), .B1(n33292), .Y(
        n21066) );
  NAND2XL U26039 ( .A(n26083), .B(n26089), .Y(n22022) );
  AOI22XL U26040 ( .A0(n21736), .A1(n22022), .B0(n26080), .B1(n21753), .Y(
        n21068) );
  OAI21XL U26041 ( .A0(n26088), .A1(n26621), .B0(n21068), .Y(n21076) );
  AOI22XL U26042 ( .A0(conv_2[223]), .A1(n21762), .B0(conv_2[238]), .B1(n21764), .Y(n21074) );
  AOI22XL U26043 ( .A0(conv_2[433]), .A1(n21765), .B0(n21751), .B1(n22012), 
        .Y(n21073) );
  AOI2BB2XL U26044 ( .B0(conv_2[403]), .B1(n21749), .A0N(n21237), .A1N(n26087), 
        .Y(n21072) );
  AOI22XL U26045 ( .A0(n22347), .A1(conv_2[298]), .B0(n16716), .B1(conv_2[313]), .Y(n21070) );
  AOI22XL U26046 ( .A0(n22759), .A1(conv_2[283]), .B0(n16673), .B1(conv_2[328]), .Y(n21069) );
  NAND2XL U26047 ( .A(n21070), .B(n21069), .Y(n26090) );
  AOI22XL U26048 ( .A0(conv_2[418]), .A1(n21763), .B0(n16663), .B1(n26090), 
        .Y(n21071) );
  NAND4XL U26049 ( .A(n21074), .B(n21073), .C(n21072), .D(n21071), .Y(n21075)
         );
  AOI211XL U26050 ( .A0(n18463), .A1(n26093), .B0(n21076), .C0(n21075), .Y(
        n21077) );
  NAND4XL U26051 ( .A(n21080), .B(n21079), .C(n21078), .D(n21077), .Y(n21083)
         );
  NAND4XL U26052 ( .A(n21082), .B(n21081), .C(n21084), .D(n21083), .Y(n21086)
         );
  NOR3XL U26053 ( .A(pool[69]), .B(n21084), .C(n21083), .Y(n21085) );
  NAND2XL U26054 ( .A(n34890), .B(pool[65]), .Y(n21090) );
  OAI21XL U26055 ( .A0(n21091), .A1(n34890), .B0(n21090), .Y(N29281) );
  ADDFX1 U26056 ( .A(DP_OP_5168J1_124_9881_n22), .B(DP_OP_5168J1_124_9881_n27), 
        .CI(n21092), .CO(n22249), .S(n20716) );
  AOI22XL U26057 ( .A0(n33563), .A1(n21093), .B0(affine_1[7]), .B1(n22250), 
        .Y(n21094) );
  NAND2XL U26058 ( .A(n21094), .B(n33077), .Y(n16506) );
  INVXL U26059 ( .A(conv_3[29]), .Y(n31309) );
  INVXL U26060 ( .A(conv_3[16]), .Y(n21110) );
  INVXL U26061 ( .A(n22846), .Y(n22209) );
  OAI22XL U26062 ( .A0(n22401), .A1(n18208), .B0(n22209), .B1(n35239), .Y(
        n21096) );
  AOI22XL U26063 ( .A0(n22370), .A1(n22402), .B0(n21100), .B1(n22396), .Y(
        n21099) );
  AOI22XL U26064 ( .A0(n22362), .A1(n22203), .B0(n22369), .B1(n22201), .Y(
        n21098) );
  AOI22XL U26065 ( .A0(n22362), .A1(n22211), .B0(n22369), .B1(n22210), .Y(
        n21101) );
  NAND3XL U26066 ( .A(conv_3[15]), .B(n34721), .C(n29678), .Y(n29427) );
  INVXL U26067 ( .A(n29427), .Y(n34720) );
  AOI32XL U26068 ( .A0(n34721), .A1(n29680), .A2(n29427), .B0(n34720), .B1(
        n30536), .Y(n21108) );
  OAI2BB1XL U26069 ( .A0N(n21108), .A1N(n21110), .B0(n21107), .Y(n21109) );
  OAI211XL U26070 ( .A0(n35576), .A1(n21110), .B0(n21109), .C0(n33550), .Y(
        n15886) );
  AOI22XL U26071 ( .A0(n21763), .A1(conv_3[405]), .B0(n21761), .B1(n34951), 
        .Y(n21122) );
  OAI2BB2XL U26072 ( .B0(n22227), .B1(n21711), .A0N(conv_3[435]), .A1N(n21752), 
        .Y(n21121) );
  AOI22XL U26073 ( .A0(conv_3[390]), .A1(n21749), .B0(conv_3[0]), .B1(n21748), 
        .Y(n21112) );
  AOI22XL U26074 ( .A0(n28559), .A1(n34962), .B0(n21756), .B1(n34964), .Y(
        n21111) );
  OAI211XL U26075 ( .A0(n21113), .A1(n21759), .B0(n21112), .C0(n21111), .Y(
        n21120) );
  AOI22XL U26076 ( .A0(conv_3[420]), .A1(n21765), .B0(n26260), .B1(n21114), 
        .Y(n21118) );
  AOI22XL U26077 ( .A0(conv_3[15]), .A1(n21766), .B0(n21464), .B1(n22235), .Y(
        n21117) );
  AOI22XL U26078 ( .A0(n28366), .A1(n34965), .B0(n16663), .B1(n34960), .Y(
        n21116) );
  NAND4XL U26079 ( .A(n21118), .B(n21117), .C(n21116), .D(n21115), .Y(n21119)
         );
  INVXL U26080 ( .A(conv_3[423]), .Y(n29688) );
  OAI22XL U26081 ( .A0(n29674), .A1(n21710), .B0(n29688), .B1(n21567), .Y(
        n21143) );
  INVXL U26082 ( .A(conv_3[18]), .Y(n29981) );
  OAI22XL U26083 ( .A0(n21123), .A1(n21712), .B0(n21729), .B1(n29981), .Y(
        n21142) );
  AOI22XL U26084 ( .A0(conv_3[438]), .A1(n21752), .B0(conv_3[408]), .B1(n21763), .Y(n21129) );
  AOI22XL U26085 ( .A0(conv_3[393]), .A1(n21749), .B0(n21761), .B1(n21124), 
        .Y(n21128) );
  AOI22XL U26086 ( .A0(n16665), .A1(n21126), .B0(n21756), .B1(n21125), .Y(
        n21127) );
  NAND3XL U26087 ( .A(n21129), .B(n21128), .C(n21127), .Y(n21141) );
  AOI22XL U26088 ( .A0(conv_3[213]), .A1(n21762), .B0(conv_3[3]), .B1(n21748), 
        .Y(n21139) );
  AOI22XL U26089 ( .A0(n22847), .A1(n21131), .B0(n21678), .B1(n21130), .Y(
        n21138) );
  AOI22XL U26090 ( .A0(n16663), .A1(n21133), .B0(n21132), .B1(n21736), .Y(
        n21137) );
  AOI22XL U26091 ( .A0(n28366), .A1(n21135), .B0(n18463), .B1(n21134), .Y(
        n21136) );
  NAND4XL U26092 ( .A(n21139), .B(n21138), .C(n21137), .D(n21136), .Y(n21140)
         );
  AOI22XL U26093 ( .A0(conv_3[406]), .A1(n21763), .B0(n21761), .B1(n21144), 
        .Y(n21146) );
  AOI22XL U26094 ( .A0(conv_3[421]), .A1(n21765), .B0(conv_3[16]), .B1(n21766), 
        .Y(n21145) );
  NAND2XL U26095 ( .A(n21146), .B(n21145), .Y(n21166) );
  INVXL U26096 ( .A(conv_3[436]), .Y(n31033) );
  OAI22XL U26097 ( .A0(n21147), .A1(n21711), .B0(n31033), .B1(n17171), .Y(
        n21165) );
  AOI22XL U26098 ( .A0(conv_3[391]), .A1(n21749), .B0(n26260), .B1(n21149), 
        .Y(n21153) );
  AOI22XL U26099 ( .A0(n28366), .A1(n21151), .B0(n21150), .B1(n21753), .Y(
        n21152) );
  NAND2XL U26100 ( .A(n21153), .B(n21152), .Y(n21164) );
  AOI22XL U26101 ( .A0(conv_3[226]), .A1(n21764), .B0(conv_3[211]), .B1(n21762), .Y(n21162) );
  AOI22XL U26102 ( .A0(n16665), .A1(n21154), .B0(conv_3[1]), .B1(n21748), .Y(
        n21161) );
  AOI22XL U26103 ( .A0(n21756), .A1(n21156), .B0(n21736), .B1(n21155), .Y(
        n21160) );
  AOI22XL U26104 ( .A0(n28559), .A1(n21158), .B0(n16663), .B1(n21157), .Y(
        n21159) );
  NAND4XL U26105 ( .A(n21162), .B(n21161), .C(n21160), .D(n21159), .Y(n21163)
         );
  AOI222XL U26106 ( .A0(n21457), .A1(pool[111]), .B0(n21457), .B1(n35011), 
        .C0(pool[111]), .C1(n35011), .Y(n21188) );
  AOI22XL U26107 ( .A0(n26260), .A1(n21167), .B0(conv_3[212]), .B1(n21762), 
        .Y(n21187) );
  AOI22XL U26108 ( .A0(conv_3[437]), .A1(n21752), .B0(conv_3[17]), .B1(n21766), 
        .Y(n21186) );
  AOI22XL U26109 ( .A0(n16665), .A1(n21169), .B0(n21756), .B1(n21168), .Y(
        n21185) );
  AOI22XL U26110 ( .A0(conv_3[407]), .A1(n21763), .B0(n21736), .B1(n21170), 
        .Y(n21171) );
  OAI21XL U26111 ( .A0(n21172), .A1(n21237), .B0(n21171), .Y(n21183) );
  AOI22XL U26112 ( .A0(n22847), .A1(n21173), .B0(conv_3[227]), .B1(n21764), 
        .Y(n21181) );
  AOI22XL U26113 ( .A0(conv_3[422]), .A1(n21765), .B0(conv_3[2]), .B1(n21748), 
        .Y(n21180) );
  AOI22XL U26114 ( .A0(n28366), .A1(n21175), .B0(n21174), .B1(n21753), .Y(
        n21179) );
  AOI22XL U26115 ( .A0(n28559), .A1(n21177), .B0(n16663), .B1(n21176), .Y(
        n21178) );
  NAND4XL U26116 ( .A(n21181), .B(n21180), .C(n21179), .D(n21178), .Y(n21182)
         );
  INVXL U26117 ( .A(pool[112]), .Y(n35013) );
  AOI222XL U26118 ( .A0(n21188), .A1(n35012), .B0(n21188), .B1(n35013), .C0(
        n35012), .C1(n35013), .Y(n21189) );
  AOI222XL U26119 ( .A0(pool[113]), .A1(n35016), .B0(pool[113]), .B1(n21189), 
        .C0(n35016), .C1(n21189), .Y(n21380) );
  INVXL U26120 ( .A(pool[114]), .Y(n22108) );
  AOI22XL U26121 ( .A0(n22847), .A1(n21191), .B0(n16663), .B1(n21190), .Y(
        n21210) );
  OAI22XL U26122 ( .A0(n21193), .A1(n21704), .B0(n21192), .B1(n16672), .Y(
        n21209) );
  AOI22XL U26123 ( .A0(conv_3[409]), .A1(n21763), .B0(n21751), .B1(n21194), 
        .Y(n21200) );
  AOI22XL U26124 ( .A0(conv_3[4]), .A1(n21748), .B0(n21678), .B1(n21195), .Y(
        n21199) );
  AOI22XL U26125 ( .A0(n16665), .A1(n21197), .B0(n28366), .B1(n21196), .Y(
        n21198) );
  NAND3XL U26126 ( .A(n21200), .B(n21199), .C(n21198), .Y(n21208) );
  AOI22XL U26127 ( .A0(conv_3[439]), .A1(n21752), .B0(conv_3[424]), .B1(n21765), .Y(n21206) );
  AOI22XL U26128 ( .A0(conv_3[229]), .A1(n21764), .B0(conv_3[19]), .B1(n21766), 
        .Y(n21205) );
  AOI22XL U26129 ( .A0(conv_3[214]), .A1(n21762), .B0(conv_3[394]), .B1(n21749), .Y(n21204) );
  AOI22XL U26130 ( .A0(n21736), .A1(n21202), .B0(n21761), .B1(n21201), .Y(
        n21203) );
  NAND4XL U26131 ( .A(n21206), .B(n21205), .C(n21204), .D(n21203), .Y(n21207)
         );
  INVXL U26132 ( .A(n22107), .Y(n21281) );
  AOI22XL U26133 ( .A0(n16663), .A1(n21212), .B0(n21756), .B1(n21211), .Y(
        n21233) );
  AOI22XL U26134 ( .A0(conv_3[217]), .A1(n21762), .B0(n21751), .B1(n21213), 
        .Y(n21215) );
  AOI22XL U26135 ( .A0(conv_3[442]), .A1(n21752), .B0(conv_3[427]), .B1(n21765), .Y(n21214) );
  OAI211XL U26136 ( .A0(n21216), .A1(n21759), .B0(n21215), .C0(n21214), .Y(
        n21224) );
  AOI22XL U26137 ( .A0(conv_3[412]), .A1(n21763), .B0(n21761), .B1(n21217), 
        .Y(n21222) );
  AOI22XL U26138 ( .A0(conv_3[397]), .A1(n21749), .B0(n21678), .B1(n21228), 
        .Y(n21221) );
  AOI22XL U26139 ( .A0(conv_3[232]), .A1(n21764), .B0(conv_3[22]), .B1(n21766), 
        .Y(n21220) );
  AOI22XL U26140 ( .A0(n28366), .A1(n21218), .B0(conv_3[7]), .B1(n21748), .Y(
        n21219) );
  NAND4XL U26141 ( .A(n21222), .B(n21221), .C(n21220), .D(n21219), .Y(n21223)
         );
  AOI211XL U26142 ( .A0(n16670), .A1(n21225), .B0(n21224), .C0(n21223), .Y(
        n21232) );
  OR2XL U26143 ( .A(n21226), .B(n36246), .Y(n21227) );
  OAI211XL U26144 ( .A0(n22743), .A1(n21228), .B0(n22847), .C0(n21227), .Y(
        n21231) );
  NAND2XL U26145 ( .A(n18463), .B(n21229), .Y(n21230) );
  NAND4XL U26146 ( .A(n21233), .B(n21232), .C(n21231), .D(n21230), .Y(n21280)
         );
  AOI22XL U26147 ( .A0(conv_3[395]), .A1(n21749), .B0(conv_3[5]), .B1(n21748), 
        .Y(n21234) );
  OAI2BB1XL U26148 ( .A0N(n21235), .A1N(n21753), .B0(n21234), .Y(n21255) );
  INVXL U26149 ( .A(conv_3[425]), .Y(n32579) );
  OAI22XL U26150 ( .A0(n21236), .A1(n21712), .B0(n32579), .B1(n21567), .Y(
        n21240) );
  INVXL U26151 ( .A(conv_3[440]), .Y(n31931) );
  OAI22XL U26152 ( .A0(n21238), .A1(n21237), .B0(n31931), .B1(n17171), .Y(
        n21239) );
  AOI211XL U26153 ( .A0(n18463), .A1(n21241), .B0(n21240), .C0(n21239), .Y(
        n21252) );
  INVXL U26154 ( .A(conv_3[410]), .Y(n32630) );
  OAI22XL U26155 ( .A0(n21242), .A1(n21711), .B0(n32630), .B1(n21536), .Y(
        n21250) );
  INVXL U26156 ( .A(conv_3[20]), .Y(n33005) );
  OAI22XL U26157 ( .A0(n28830), .A1(n21556), .B0(n33005), .B1(n21729), .Y(
        n21249) );
  OAI22XL U26158 ( .A0(n21244), .A1(n28553), .B0(n21243), .B1(n28349), .Y(
        n21248) );
  OAI22XL U26159 ( .A0(n21246), .A1(n21759), .B0(n21245), .B1(n26621), .Y(
        n21247) );
  NOR4XL U26160 ( .A(n21250), .B(n21249), .C(n21248), .D(n21247), .Y(n21251)
         );
  OAI211XL U26161 ( .A0(n21253), .A1(n21704), .B0(n21252), .C0(n21251), .Y(
        n21254) );
  AOI211XL U26162 ( .A0(conv_3[230]), .A1(n21764), .B0(n21255), .C0(n21254), 
        .Y(n21256) );
  INVXL U26163 ( .A(n21256), .Y(n21375) );
  AOI22XL U26164 ( .A0(n28366), .A1(n21258), .B0(n16663), .B1(n21257), .Y(
        n21261) );
  NAND2XL U26165 ( .A(n21756), .B(n21259), .Y(n21260) );
  OAI211XL U26166 ( .A0(n21262), .A1(n21759), .B0(n21261), .C0(n21260), .Y(
        n21279) );
  NAND2XL U26167 ( .A(n22713), .B(n21263), .Y(n21264) );
  OAI22XL U26168 ( .A0(n28277), .A1(n21264), .B0(n32093), .B1(n21710), .Y(
        n21278) );
  AOI22XL U26169 ( .A0(conv_3[216]), .A1(n21762), .B0(conv_3[411]), .B1(n21763), .Y(n21268) );
  AOI22XL U26170 ( .A0(n16665), .A1(n21266), .B0(n21265), .B1(n21753), .Y(
        n21267) );
  NAND2XL U26171 ( .A(n21268), .B(n21267), .Y(n21277) );
  AOI22XL U26172 ( .A0(conv_3[396]), .A1(n21749), .B0(n21751), .B1(n21269), 
        .Y(n21275) );
  AOI22XL U26173 ( .A0(n21748), .A1(conv_3[6]), .B0(n21761), .B1(n21270), .Y(
        n21274) );
  AOI22XL U26174 ( .A0(conv_3[441]), .A1(n21752), .B0(conv_3[21]), .B1(n21766), 
        .Y(n21273) );
  AOI22XL U26175 ( .A0(n28559), .A1(n21271), .B0(conv_3[426]), .B1(n21765), 
        .Y(n21272) );
  NAND4XL U26176 ( .A(n21275), .B(n21274), .C(n21273), .D(n21272), .Y(n21276)
         );
  AOI22XL U26177 ( .A0(conv_3[219]), .A1(n21762), .B0(conv_3[9]), .B1(n21748), 
        .Y(n21284) );
  AOI22XL U26178 ( .A0(conv_3[444]), .A1(n21752), .B0(n21761), .B1(n21282), 
        .Y(n21283) );
  OAI211XL U26179 ( .A0(n21285), .A1(n21704), .B0(n21284), .C0(n21283), .Y(
        n21303) );
  AOI22XL U26180 ( .A0(conv_3[24]), .A1(n21766), .B0(n21751), .B1(n21286), .Y(
        n21301) );
  AOI22XL U26181 ( .A0(n16665), .A1(n21288), .B0(n16663), .B1(n21287), .Y(
        n21294) );
  OAI22XL U26182 ( .A0(n30694), .A1(n21710), .B0(n32555), .B1(n21536), .Y(
        n21293) );
  INVXL U26183 ( .A(conv_3[429]), .Y(n35777) );
  OAI22XL U26184 ( .A0(n35777), .A1(n21567), .B0(n32047), .B1(n21731), .Y(
        n21292) );
  OAI22XL U26185 ( .A0(n21290), .A1(n16672), .B0(n21289), .B1(n21759), .Y(
        n21291) );
  NOR4BXL U26186 ( .AN(n21294), .B(n21293), .C(n21292), .D(n21291), .Y(n21300)
         );
  OAI22XL U26187 ( .A0(n21678), .A1(n21298), .B0(n21358), .B1(n21297), .Y(
        n21299) );
  NAND3XL U26188 ( .A(n21301), .B(n21300), .C(n21299), .Y(n21302) );
  AOI211XL U26189 ( .A0(n28366), .A1(n21304), .B0(n21303), .C0(n21302), .Y(
        n21447) );
  AOI22XL U26190 ( .A0(n16663), .A1(n21306), .B0(n21736), .B1(n21305), .Y(
        n21309) );
  NAND2XL U26191 ( .A(n18463), .B(n21307), .Y(n21308) );
  OAI211XL U26192 ( .A0(n21310), .A1(n21704), .B0(n21309), .C0(n21308), .Y(
        n21328) );
  OAI22XL U26193 ( .A0(n21313), .A1(n21711), .B0(n21312), .B1(n21311), .Y(
        n21327) );
  AOI22XL U26194 ( .A0(conv_3[446]), .A1(n21752), .B0(n21761), .B1(n21314), 
        .Y(n21316) );
  AOI22XL U26195 ( .A0(conv_3[236]), .A1(n21764), .B0(conv_3[11]), .B1(n21748), 
        .Y(n21315) );
  OAI211XL U26196 ( .A0(n21317), .A1(n28553), .B0(n21316), .C0(n21315), .Y(
        n21326) );
  AOI22XL U26197 ( .A0(conv_3[416]), .A1(n21763), .B0(conv_3[401]), .B1(n21749), .Y(n21324) );
  AOI22XL U26198 ( .A0(conv_3[221]), .A1(n21762), .B0(n21678), .B1(n21318), 
        .Y(n21323) );
  AOI22XL U26199 ( .A0(conv_3[431]), .A1(n21765), .B0(conv_3[26]), .B1(n21766), 
        .Y(n21322) );
  AOI22XL U26200 ( .A0(n28366), .A1(n21320), .B0(n26260), .B1(n21319), .Y(
        n21321) );
  NAND4XL U26201 ( .A(n21324), .B(n21323), .C(n21322), .D(n21321), .Y(n21325)
         );
  NOR4XL U26202 ( .A(n21328), .B(n21327), .C(n21326), .D(n21325), .Y(n21450)
         );
  AOI22XL U26203 ( .A0(conv_3[233]), .A1(n21764), .B0(n26260), .B1(n21329), 
        .Y(n21330) );
  OAI2BB1XL U26204 ( .A0N(n22847), .A1N(n21331), .B0(n21330), .Y(n21332) );
  AOI22XL U26205 ( .A0(conv_3[428]), .A1(n21765), .B0(conv_3[23]), .B1(n21766), 
        .Y(n21349) );
  AOI22XL U26206 ( .A0(conv_3[413]), .A1(n21763), .B0(conv_3[8]), .B1(n21748), 
        .Y(n21348) );
  AOI22XL U26207 ( .A0(n16665), .A1(n21335), .B0(n21756), .B1(n21334), .Y(
        n21338) );
  NAND2XL U26208 ( .A(n28324), .B(n21336), .Y(n21337) );
  OAI211XL U26209 ( .A0(n21339), .A1(n28349), .B0(n21338), .C0(n21337), .Y(
        n21345) );
  AOI22XL U26210 ( .A0(conv_3[218]), .A1(n21762), .B0(conv_3[398]), .B1(n21749), .Y(n21342) );
  AOI22XL U26211 ( .A0(conv_3[443]), .A1(n21752), .B0(n21761), .B1(n21340), 
        .Y(n21341) );
  OAI211XL U26212 ( .A0(n21343), .A1(n21759), .B0(n21342), .C0(n21341), .Y(
        n21344) );
  AOI211XL U26213 ( .A0(n18463), .A1(n21346), .B0(n21345), .C0(n21344), .Y(
        n21347) );
  NAND4XL U26214 ( .A(n21350), .B(n21349), .C(n21348), .D(n21347), .Y(n21445)
         );
  INVXL U26215 ( .A(conv_3[445]), .Y(n33763) );
  OAI22XL U26216 ( .A0(n33763), .A1(n17171), .B0(n31256), .B1(n21729), .Y(
        n21351) );
  AOI2BB1XL U26217 ( .A0N(n21352), .A1N(n21704), .B0(n21351), .Y(n21373) );
  AOI22XL U26218 ( .A0(conv_3[415]), .A1(n21763), .B0(n21761), .B1(n21353), 
        .Y(n21355) );
  AOI22XL U26219 ( .A0(conv_3[430]), .A1(n21765), .B0(conv_3[220]), .B1(n21762), .Y(n21354) );
  OAI211XL U26220 ( .A0(n21356), .A1(n26621), .B0(n21355), .C0(n21354), .Y(
        n21370) );
  AOI2BB2XL U26221 ( .B0(n21748), .B1(conv_3[10]), .A0N(n21357), .A1N(n21711), 
        .Y(n21368) );
  AOI22XL U26222 ( .A0(conv_3[400]), .A1(n21749), .B0(n26260), .B1(n21360), 
        .Y(n21367) );
  AOI22XL U26223 ( .A0(n18463), .A1(n21362), .B0(n16663), .B1(n21361), .Y(
        n21366) );
  AOI22XL U26224 ( .A0(n16665), .A1(n21364), .B0(n21736), .B1(n21363), .Y(
        n21365) );
  NAND4XL U26225 ( .A(n21368), .B(n21367), .C(n21366), .D(n21365), .Y(n21369)
         );
  AOI211XL U26226 ( .A0(n21371), .A1(n21753), .B0(n21370), .C0(n21369), .Y(
        n21372) );
  OAI211XL U26227 ( .A0(n29166), .A1(n21710), .B0(n21373), .C0(n21372), .Y(
        n21444) );
  NOR4XL U26228 ( .A(n21375), .B(n21374), .C(n21445), .D(n21444), .Y(n21376)
         );
  NAND4XL U26229 ( .A(n21377), .B(n21447), .C(n21450), .D(n21376), .Y(n21378)
         );
  AOI22XL U26230 ( .A0(conv_3[449]), .A1(n21752), .B0(n21761), .B1(n21381), 
        .Y(n21401) );
  AOI22XL U26231 ( .A0(conv_3[239]), .A1(n21764), .B0(conv_3[404]), .B1(n21749), .Y(n21400) );
  AOI22XL U26232 ( .A0(conv_3[224]), .A1(n21762), .B0(conv_3[419]), .B1(n21763), .Y(n21384) );
  AOI22XL U26233 ( .A0(n26260), .A1(n21382), .B0(conv_3[14]), .B1(n21748), .Y(
        n21383) );
  OAI211XL U26234 ( .A0(n21385), .A1(n21759), .B0(n21384), .C0(n21383), .Y(
        n21386) );
  AOI21XL U26235 ( .A0(n16663), .A1(n21387), .B0(n21386), .Y(n21399) );
  OAI22XL U26236 ( .A0(n21388), .A1(n21711), .B0(n31309), .B1(n21729), .Y(
        n21397) );
  INVXL U26237 ( .A(conv_3[434]), .Y(n32162) );
  OAI22XL U26238 ( .A0(n21389), .A1(n26621), .B0(n32162), .B1(n21567), .Y(
        n21396) );
  INVXL U26239 ( .A(n21753), .Y(n21703) );
  OAI22XL U26240 ( .A0(n21391), .A1(n21703), .B0(n21390), .B1(n28553), .Y(
        n21395) );
  OAI2BB2XL U26241 ( .B0(n21393), .B1(n21704), .A0N(n18463), .A1N(n21392), .Y(
        n21394) );
  NOR4XL U26242 ( .A(n21397), .B(n21396), .C(n21395), .D(n21394), .Y(n21398)
         );
  NAND4XL U26243 ( .A(n21401), .B(n21400), .C(n21399), .D(n21398), .Y(n21453)
         );
  AOI22XL U26244 ( .A0(conv_3[403]), .A1(n21749), .B0(n21761), .B1(n21402), 
        .Y(n21422) );
  AOI22XL U26245 ( .A0(conv_3[223]), .A1(n21762), .B0(n21751), .B1(n21403), 
        .Y(n21421) );
  AOI22XL U26246 ( .A0(n16665), .A1(n21405), .B0(n28366), .B1(n21404), .Y(
        n21420) );
  AOI22XL U26247 ( .A0(conv_3[238]), .A1(n21764), .B0(conv_3[28]), .B1(n21766), 
        .Y(n21406) );
  OAI21XL U26248 ( .A0(n21407), .A1(n21704), .B0(n21406), .Y(n21417) );
  AOI22XL U26249 ( .A0(conv_3[448]), .A1(n21752), .B0(conv_3[13]), .B1(n21748), 
        .Y(n21415) );
  AOI22XL U26250 ( .A0(conv_3[433]), .A1(n21765), .B0(conv_3[418]), .B1(n21763), .Y(n21414) );
  AOI2BB2XL U26251 ( .B0(n21736), .B1(n21409), .A0N(n21408), .A1N(n16672), .Y(
        n21413) );
  AOI22XL U26252 ( .A0(n16663), .A1(n21411), .B0(n21410), .B1(n21753), .Y(
        n21412) );
  NAND4XL U26253 ( .A(n21415), .B(n21414), .C(n21413), .D(n21412), .Y(n21416)
         );
  AOI211XL U26254 ( .A0(n22847), .A1(n21418), .B0(n21417), .C0(n21416), .Y(
        n21419) );
  NAND4XL U26255 ( .A(n21422), .B(n21421), .C(n21420), .D(n21419), .Y(n21448)
         );
  AOI22XL U26256 ( .A0(conv_3[447]), .A1(n21752), .B0(n21761), .B1(n21423), 
        .Y(n21443) );
  AOI22XL U26257 ( .A0(conv_3[222]), .A1(n21762), .B0(n21725), .B1(n21424), 
        .Y(n21442) );
  AOI22XL U26258 ( .A0(conv_3[237]), .A1(n21764), .B0(conv_3[27]), .B1(n21766), 
        .Y(n21427) );
  AOI22XL U26259 ( .A0(conv_3[417]), .A1(n21763), .B0(n26260), .B1(n21425), 
        .Y(n21426) );
  OAI211XL U26260 ( .A0(n21428), .A1(n26621), .B0(n21427), .C0(n21426), .Y(
        n21429) );
  AOI2BB1XL U26261 ( .A0N(n21430), .A1N(n28553), .B0(n21429), .Y(n21441) );
  AOI22XL U26262 ( .A0(n28559), .A1(n21432), .B0(n21431), .B1(n21753), .Y(
        n21439) );
  INVXL U26263 ( .A(conv_3[432]), .Y(n32586) );
  INVXL U26264 ( .A(conv_3[12]), .Y(n28640) );
  OAI22XL U26265 ( .A0(n32586), .A1(n21567), .B0(n28640), .B1(n21730), .Y(
        n21438) );
  INVXL U26266 ( .A(conv_3[402]), .Y(n33698) );
  OAI22XL U26267 ( .A0(n21433), .A1(n21704), .B0(n33698), .B1(n21731), .Y(
        n21437) );
  OAI22XL U26268 ( .A0(n21435), .A1(n21759), .B0(n21434), .B1(n28349), .Y(
        n21436) );
  NOR4BXL U26269 ( .AN(n21439), .B(n21438), .C(n21437), .D(n21436), .Y(n21440)
         );
  NAND4XL U26270 ( .A(n21443), .B(n21442), .C(n21441), .D(n21440), .Y(n21446)
         );
  NOR3XL U26271 ( .A(pool[114]), .B(n21448), .C(n21446), .Y(n21452) );
  NAND4BXL U26272 ( .AN(n21447), .B(n21446), .C(n21445), .D(n21444), .Y(n21449) );
  NAND4BBXL U26273 ( .AN(n21450), .BN(n21449), .C(pool[114]), .D(n21448), .Y(
        n21451) );
  NAND2XL U26274 ( .A(n35014), .B(pool[110]), .Y(n21456) );
  OAI21XL U26275 ( .A0(n21457), .A1(n35014), .B0(n21456), .Y(N29326) );
  INVXL U26276 ( .A(conv_1[405]), .Y(n33522) );
  INVXL U26277 ( .A(conv_1[0]), .Y(n26959) );
  OAI22XL U26278 ( .A0(n33522), .A1(n21536), .B0(n26959), .B1(n21730), .Y(
        n21477) );
  INVXL U26279 ( .A(conv_1[390]), .Y(n30651) );
  OAI22XL U26280 ( .A0(n25305), .A1(n21711), .B0(n21731), .B1(n30651), .Y(
        n21476) );
  AOI22XL U26281 ( .A0(n21765), .A1(conv_1[420]), .B0(n21761), .B1(n25297), 
        .Y(n21462) );
  AOI22XL U26282 ( .A0(n16665), .A1(n21460), .B0(n16663), .B1(n21459), .Y(
        n21461) );
  OAI211XL U26283 ( .A0(n21463), .A1(n21704), .B0(n21462), .C0(n21461), .Y(
        n21475) );
  AOI22XL U26284 ( .A0(conv_1[435]), .A1(n21752), .B0(n21464), .B1(n25298), 
        .Y(n21473) );
  AOI22XL U26285 ( .A0(conv_1[15]), .A1(n21766), .B0(n21751), .B1(n21465), .Y(
        n21472) );
  AOI2BB2XL U26286 ( .B0(n18463), .B1(n21467), .A0N(n21466), .A1N(n28575), .Y(
        n21471) );
  AOI22XL U26287 ( .A0(n28366), .A1(n21469), .B0(n21468), .B1(n21736), .Y(
        n21470) );
  NAND4XL U26288 ( .A(n21473), .B(n21472), .C(n21471), .D(n21470), .Y(n21474)
         );
  AOI22XL U26289 ( .A0(conv_1[408]), .A1(n21763), .B0(conv_1[213]), .B1(n21762), .Y(n21478) );
  OAI2BB1XL U26290 ( .A0N(n21761), .A1N(n22635), .B0(n21478), .Y(n21495) );
  AOI22XL U26291 ( .A0(n22847), .A1(n21479), .B0(conv_1[228]), .B1(n21764), 
        .Y(n21493) );
  AOI22XL U26292 ( .A0(conv_1[393]), .A1(n21749), .B0(conv_1[3]), .B1(n21748), 
        .Y(n21492) );
  AOI22XL U26293 ( .A0(n28559), .A1(n21480), .B0(n22638), .B1(n21753), .Y(
        n21491) );
  AOI22XL U26294 ( .A0(conv_1[438]), .A1(n21752), .B0(n21751), .B1(n22643), 
        .Y(n21489) );
  AOI22XL U26295 ( .A0(conv_1[423]), .A1(n21765), .B0(n21756), .B1(n21481), 
        .Y(n21488) );
  AOI22XL U26296 ( .A0(n16665), .A1(n21483), .B0(n28366), .B1(n21482), .Y(
        n21487) );
  AOI22XL U26297 ( .A0(n21736), .A1(n21485), .B0(n16663), .B1(n21484), .Y(
        n21486) );
  NAND4XL U26298 ( .A(n21493), .B(n21492), .C(n21491), .D(n21490), .Y(n21494)
         );
  INVXL U26299 ( .A(conv_1[391]), .Y(n30671) );
  OAI22XL U26300 ( .A0(n18196), .A1(n21496), .B0(n30671), .B1(n21731), .Y(
        n21514) );
  INVXL U26301 ( .A(conv_1[226]), .Y(n23953) );
  OAI22XL U26302 ( .A0(n21497), .A1(n16672), .B0(n23953), .B1(n21710), .Y(
        n21513) );
  INVXL U26303 ( .A(conv_1[1]), .Y(n27433) );
  OAI22XL U26304 ( .A0(n22683), .A1(n21711), .B0(n21730), .B1(n27433), .Y(
        n21500) );
  INVXL U26305 ( .A(conv_1[16]), .Y(n27465) );
  OAI22XL U26306 ( .A0(n27465), .A1(n21729), .B0(n26285), .B1(n21498), .Y(
        n21499) );
  AOI211XL U26307 ( .A0(n21736), .A1(n21501), .B0(n21500), .C0(n21499), .Y(
        n21502) );
  OAI21XL U26308 ( .A0(n21503), .A1(n26621), .B0(n21502), .Y(n21512) );
  AOI22XL U26309 ( .A0(conv_1[406]), .A1(n21763), .B0(conv_1[211]), .B1(n21762), .Y(n21510) );
  AOI22XL U26310 ( .A0(conv_1[436]), .A1(n21752), .B0(conv_1[421]), .B1(n21765), .Y(n21509) );
  AOI2BB2XL U26311 ( .B0(n22696), .B1(n21753), .A0N(n21504), .A1N(n28553), .Y(
        n21508) );
  AOI22XL U26312 ( .A0(n16663), .A1(n21506), .B0(n21756), .B1(n21505), .Y(
        n21507) );
  NAND4XL U26313 ( .A(n21510), .B(n21509), .C(n21508), .D(n21507), .Y(n21511)
         );
  AOI222XL U26314 ( .A0(pool[21]), .A1(n21793), .B0(pool[21]), .B1(n34812), 
        .C0(n21793), .C1(n34812), .Y(n21533) );
  AOI22XL U26315 ( .A0(conv_1[227]), .A1(n21764), .B0(conv_1[212]), .B1(n21762), .Y(n21532) );
  AOI22XL U26316 ( .A0(conv_1[392]), .A1(n21749), .B0(conv_1[2]), .B1(n21748), 
        .Y(n21531) );
  AOI22XL U26317 ( .A0(n28559), .A1(n21516), .B0(n21756), .B1(n21515), .Y(
        n21530) );
  AOI22XL U26318 ( .A0(conv_1[407]), .A1(n21763), .B0(n26260), .B1(n21517), 
        .Y(n21518) );
  OAI2BB1XL U26319 ( .A0N(n21725), .A1N(n22657), .B0(n21518), .Y(n21528) );
  AOI22XL U26320 ( .A0(conv_1[437]), .A1(n21752), .B0(conv_1[422]), .B1(n21765), .Y(n21526) );
  AOI22XL U26321 ( .A0(n28366), .A1(n21519), .B0(n21761), .B1(n22662), .Y(
        n21525) );
  AOI22XL U26322 ( .A0(n16663), .A1(n21521), .B0(n21736), .B1(n21520), .Y(
        n21524) );
  AOI22XL U26323 ( .A0(n16665), .A1(n21522), .B0(n22655), .B1(n21753), .Y(
        n21523) );
  NAND4XL U26324 ( .A(n21526), .B(n21525), .C(n21524), .D(n21523), .Y(n21527)
         );
  AOI211XL U26325 ( .A0(conv_1[17]), .A1(n21766), .B0(n21528), .C0(n21527), 
        .Y(n21529) );
  NAND4XL U26326 ( .A(n21532), .B(n21531), .C(n21530), .D(n21529), .Y(n34814)
         );
  AOI222XL U26327 ( .A0(n21533), .A1(n34814), .B0(n21533), .B1(n34816), .C0(
        n34814), .C1(n34816), .Y(n21534) );
  AOI222XL U26328 ( .A0(pool[23]), .A1(n22098), .B0(pool[23]), .B1(n21534), 
        .C0(n22098), .C1(n21534), .Y(n21702) );
  OAI22XL U26329 ( .A0(n35486), .A1(n21536), .B0(n26285), .B1(n21535), .Y(
        n21555) );
  INVXL U26330 ( .A(conv_1[229]), .Y(n23914) );
  OAI22XL U26331 ( .A0(n22498), .A1(n21703), .B0(n23914), .B1(n21710), .Y(
        n21554) );
  OAI2BB2XL U26332 ( .B0(n27455), .B1(n21729), .A0N(conv_1[4]), .A1N(n21748), 
        .Y(n21540) );
  OAI22XL U26333 ( .A0(n28277), .A1(n21538), .B0(n18196), .B1(n21537), .Y(
        n21539) );
  AOI211XL U26334 ( .A0(n28324), .A1(n21541), .B0(n21540), .C0(n21539), .Y(
        n21542) );
  OAI2BB1XL U26335 ( .A0N(n18463), .A1N(n21543), .B0(n21542), .Y(n21553) );
  AOI22XL U26336 ( .A0(conv_1[394]), .A1(n21749), .B0(conv_1[439]), .B1(n21752), .Y(n21551) );
  AOI22XL U26337 ( .A0(conv_1[214]), .A1(n21762), .B0(conv_1[424]), .B1(n21765), .Y(n21550) );
  AOI22XL U26338 ( .A0(n16665), .A1(n21545), .B0(n21736), .B1(n21544), .Y(
        n21549) );
  AOI22XL U26339 ( .A0(n16663), .A1(n21547), .B0(n21756), .B1(n21546), .Y(
        n21548) );
  NAND4XL U26340 ( .A(n21551), .B(n21550), .C(n21549), .D(n21548), .Y(n21552)
         );
  NOR4XL U26341 ( .A(n21555), .B(n21554), .C(n21553), .D(n21552), .Y(n22096)
         );
  INVXL U26342 ( .A(conv_1[21]), .Y(n27349) );
  INVXL U26343 ( .A(conv_1[396]), .Y(n29273) );
  OAI22XL U26344 ( .A0(n27349), .A1(n21729), .B0(n29273), .B1(n21731), .Y(
        n21578) );
  INVXL U26345 ( .A(conv_1[216]), .Y(n23308) );
  OAI22XL U26346 ( .A0(n23308), .A1(n21556), .B0(n29267), .B1(n21710), .Y(
        n21577) );
  AOI22XL U26347 ( .A0(conv_1[441]), .A1(n21752), .B0(conv_1[6]), .B1(n21748), 
        .Y(n21559) );
  NAND2XL U26348 ( .A(n16670), .B(n21557), .Y(n21558) );
  OAI211XL U26349 ( .A0(n21564), .A1(n28575), .B0(n21559), .C0(n21558), .Y(
        n21576) );
  OAI22XL U26350 ( .A0(n21561), .A1(n21704), .B0(n21560), .B1(n16672), .Y(
        n21574) );
  AOI22XL U26351 ( .A0(n28366), .A1(n21563), .B0(n16663), .B1(n21562), .Y(
        n21573) );
  AOI22XL U26352 ( .A0(conv_1[411]), .A1(n21763), .B0(n21761), .B1(n22460), 
        .Y(n21572) );
  AOI21XL U26353 ( .A0(n21565), .A1(n21564), .B0(n28277), .Y(n21569) );
  INVXL U26354 ( .A(conv_1[426]), .Y(n35503) );
  OAI22XL U26355 ( .A0(n35503), .A1(n21567), .B0(n26285), .B1(n21566), .Y(
        n21568) );
  AOI211XL U26356 ( .A0(n21736), .A1(n21570), .B0(n21569), .C0(n21568), .Y(
        n21571) );
  NAND4BXL U26357 ( .AN(n21574), .B(n21573), .C(n21572), .D(n21571), .Y(n21575) );
  NOR4XL U26358 ( .A(n21578), .B(n21577), .C(n21576), .D(n21575), .Y(n21695)
         );
  AOI22XL U26359 ( .A0(n28324), .A1(n21580), .B0(n16663), .B1(n21579), .Y(
        n21582) );
  AOI32XL U26360 ( .A0(n21583), .A1(n21582), .A2(n21581), .B0(n28277), .B1(
        n21582), .Y(n21596) );
  AOI22XL U26361 ( .A0(conv_1[232]), .A1(n21764), .B0(conv_1[427]), .B1(n21765), .Y(n21594) );
  AOI22XL U26362 ( .A0(conv_1[412]), .A1(n21763), .B0(conv_1[217]), .B1(n21762), .Y(n21593) );
  AOI22XL U26363 ( .A0(n28559), .A1(n21585), .B0(n21736), .B1(n21584), .Y(
        n21592) );
  AOI22XL U26364 ( .A0(n21748), .A1(conv_1[7]), .B0(n21751), .B1(n22626), .Y(
        n21590) );
  AOI22XL U26365 ( .A0(conv_1[397]), .A1(n21749), .B0(n21761), .B1(n22611), 
        .Y(n21589) );
  AOI22XL U26366 ( .A0(conv_1[442]), .A1(n21752), .B0(n21678), .B1(n22623), 
        .Y(n21588) );
  AOI22XL U26367 ( .A0(conv_1[22]), .A1(n21766), .B0(n21756), .B1(n21586), .Y(
        n21587) );
  NAND4XL U26368 ( .A(n21594), .B(n21593), .C(n21592), .D(n21591), .Y(n21595)
         );
  AOI211XL U26369 ( .A0(n16665), .A1(n21597), .B0(n21596), .C0(n21595), .Y(
        n21698) );
  AOI22XL U26370 ( .A0(n28324), .A1(n21599), .B0(n16663), .B1(n21598), .Y(
        n21609) );
  AOI22XL U26371 ( .A0(n16670), .A1(n21601), .B0(n21600), .B1(n21736), .Y(
        n21608) );
  AOI22XL U26372 ( .A0(n21765), .A1(conv_1[425]), .B0(n21761), .B1(n22568), 
        .Y(n21607) );
  INVXL U26373 ( .A(n22582), .Y(n21602) );
  AOI221XL U26374 ( .A0(n21602), .A1(n36246), .B0(n22579), .B1(n21688), .C0(
        n28277), .Y(n21604) );
  INVXL U26375 ( .A(conv_1[395]), .Y(n29279) );
  OAI22XL U26376 ( .A0(n22578), .A1(n21712), .B0(n29279), .B1(n21731), .Y(
        n21603) );
  AOI211XL U26377 ( .A0(n21756), .A1(n21605), .B0(n21604), .C0(n21603), .Y(
        n21606) );
  NAND4XL U26378 ( .A(n21609), .B(n21608), .C(n21607), .D(n21606), .Y(n21616)
         );
  AOI22XL U26379 ( .A0(conv_1[20]), .A1(n21766), .B0(conv_1[230]), .B1(n21764), 
        .Y(n21614) );
  AOI22XL U26380 ( .A0(conv_1[215]), .A1(n21762), .B0(conv_1[5]), .B1(n21748), 
        .Y(n21613) );
  AOI22XL U26381 ( .A0(conv_1[440]), .A1(n21752), .B0(n21678), .B1(n22582), 
        .Y(n21612) );
  AOI22XL U26382 ( .A0(n28559), .A1(n21610), .B0(conv_1[410]), .B1(n21763), 
        .Y(n21611) );
  NAND4XL U26383 ( .A(n21614), .B(n21613), .C(n21612), .D(n21611), .Y(n21615)
         );
  NOR4XL U26384 ( .A(n22096), .B(n21695), .C(n21698), .D(n21697), .Y(n21701)
         );
  AOI22XL U26385 ( .A0(conv_1[413]), .A1(n21763), .B0(n21678), .B1(n22557), 
        .Y(n21635) );
  AOI22XL U26386 ( .A0(conv_1[23]), .A1(n21766), .B0(conv_1[398]), .B1(n21749), 
        .Y(n21634) );
  AOI221XL U26387 ( .A0(n21617), .A1(n36246), .B0(n22556), .B1(n21688), .C0(
        n28277), .Y(n21621) );
  AOI22XL U26388 ( .A0(conv_1[428]), .A1(n21765), .B0(n21761), .B1(n22560), 
        .Y(n21619) );
  NAND2XL U26389 ( .A(conv_1[8]), .B(n21748), .Y(n21618) );
  OAI211XL U26390 ( .A0(n22555), .A1(n21712), .B0(n21619), .C0(n21618), .Y(
        n21620) );
  AOI211XL U26391 ( .A0(n16670), .A1(n21622), .B0(n21621), .C0(n21620), .Y(
        n21633) );
  AOI22XL U26392 ( .A0(conv_1[218]), .A1(n21762), .B0(conv_1[233]), .B1(n21764), .Y(n21631) );
  AOI22XL U26393 ( .A0(conv_1[443]), .A1(n21752), .B0(n21623), .B1(n21736), 
        .Y(n21630) );
  AOI22XL U26394 ( .A0(n28366), .A1(n21625), .B0(n21756), .B1(n21624), .Y(
        n21629) );
  AOI22XL U26395 ( .A0(n28559), .A1(n21627), .B0(n16663), .B1(n21626), .Y(
        n21628) );
  NAND4XL U26396 ( .A(n21635), .B(n21634), .C(n21633), .D(n21632), .Y(n21781)
         );
  OAI22XL U26397 ( .A0(n21637), .A1(n21704), .B0(n21636), .B1(n26621), .Y(
        n21638) );
  AOI21XL U26398 ( .A0(n22487), .A1(n21753), .B0(n21638), .Y(n21653) );
  AOI22XL U26399 ( .A0(n22847), .A1(n21639), .B0(n21761), .B1(n22490), .Y(
        n21641) );
  AOI22XL U26400 ( .A0(conv_1[430]), .A1(n21765), .B0(conv_1[445]), .B1(n21752), .Y(n21640) );
  OAI211XL U26401 ( .A0(n21642), .A1(n21759), .B0(n21641), .C0(n21640), .Y(
        n21650) );
  AOI22XL U26402 ( .A0(conv_1[400]), .A1(n21749), .B0(n26260), .B1(n21643), 
        .Y(n21648) );
  AOI22XL U26403 ( .A0(conv_1[25]), .A1(n21766), .B0(conv_1[220]), .B1(n21762), 
        .Y(n21647) );
  AOI22XL U26404 ( .A0(conv_1[415]), .A1(n21763), .B0(conv_1[10]), .B1(n21748), 
        .Y(n21646) );
  AOI22XL U26405 ( .A0(n28559), .A1(n21644), .B0(conv_1[235]), .B1(n21764), 
        .Y(n21645) );
  NAND4XL U26406 ( .A(n21648), .B(n21647), .C(n21646), .D(n21645), .Y(n21649)
         );
  AOI211XL U26407 ( .A0(n16663), .A1(n21651), .B0(n21650), .C0(n21649), .Y(
        n21652) );
  OAI211XL U26408 ( .A0(n21654), .A1(n28553), .B0(n21653), .C0(n21652), .Y(
        n21782) );
  AOI22XL U26409 ( .A0(conv_1[399]), .A1(n21749), .B0(conv_1[429]), .B1(n21765), .Y(n21672) );
  AOI22XL U26410 ( .A0(conv_1[414]), .A1(n21763), .B0(conv_1[9]), .B1(n21748), 
        .Y(n21671) );
  AOI22XL U26411 ( .A0(conv_1[234]), .A1(n21764), .B0(n21751), .B1(n22521), 
        .Y(n21656) );
  AOI22XL U26412 ( .A0(conv_1[219]), .A1(n21762), .B0(conv_1[444]), .B1(n21752), .Y(n21655) );
  OAI211XL U26413 ( .A0(n21657), .A1(n21759), .B0(n21656), .C0(n21655), .Y(
        n21658) );
  AOI2BB1XL U26414 ( .A0N(n21659), .A1N(n16672), .B0(n21658), .Y(n21670) );
  AOI22XL U26415 ( .A0(n21678), .A1(n22525), .B0(n21761), .B1(n22532), .Y(
        n21668) );
  INVXL U26416 ( .A(conv_1[24]), .Y(n27611) );
  OAI22XL U26417 ( .A0(n21660), .A1(n28349), .B0(n27611), .B1(n21729), .Y(
        n21667) );
  OAI22XL U26418 ( .A0(n21662), .A1(n21704), .B0(n28277), .B1(n21661), .Y(
        n21666) );
  OAI22XL U26419 ( .A0(n21664), .A1(n28553), .B0(n21663), .B1(n26621), .Y(
        n21665) );
  NOR4BXL U26420 ( .AN(n21668), .B(n21667), .C(n21666), .D(n21665), .Y(n21669)
         );
  NAND4XL U26421 ( .A(n21672), .B(n21671), .C(n21670), .D(n21669), .Y(n21785)
         );
  AOI22XL U26422 ( .A0(n28366), .A1(n21674), .B0(n21756), .B1(n21673), .Y(
        n21694) );
  AOI22XL U26423 ( .A0(conv_1[221]), .A1(n21762), .B0(conv_1[416]), .B1(n21763), .Y(n21676) );
  AOI22XL U26424 ( .A0(conv_1[446]), .A1(n21752), .B0(n21751), .B1(n22595), 
        .Y(n21675) );
  OAI211XL U26425 ( .A0(n21677), .A1(n21759), .B0(n21676), .C0(n21675), .Y(
        n21685) );
  AOI22XL U26426 ( .A0(conv_1[11]), .A1(n21748), .B0(n21761), .B1(n22590), .Y(
        n21683) );
  AOI22XL U26427 ( .A0(conv_1[26]), .A1(n21766), .B0(conv_1[236]), .B1(n21764), 
        .Y(n21682) );
  AOI22XL U26428 ( .A0(conv_1[401]), .A1(n21749), .B0(n21678), .B1(n22599), 
        .Y(n21681) );
  AOI22XL U26429 ( .A0(n16665), .A1(n21679), .B0(conv_1[431]), .B1(n21765), 
        .Y(n21680) );
  NAND4XL U26430 ( .A(n21683), .B(n21682), .C(n21681), .D(n21680), .Y(n21684)
         );
  AOI211XL U26431 ( .A0(n16663), .A1(n21686), .B0(n21685), .C0(n21684), .Y(
        n21693) );
  NAND2XL U26432 ( .A(n18463), .B(n21687), .Y(n21692) );
  NAND2XL U26433 ( .A(n21689), .B(n21688), .Y(n21690) );
  OAI211XL U26434 ( .A0(n22765), .A1(n22599), .B0(n22847), .C0(n21690), .Y(
        n21691) );
  NAND4XL U26435 ( .A(n21694), .B(n21693), .C(n21692), .D(n21691), .Y(n21784)
         );
  NOR4BBXL U26436 ( .AN(n22096), .BN(n21695), .C(n21785), .D(n21784), .Y(
        n21696) );
  NAND4XL U26437 ( .A(n21699), .B(n21698), .C(n21697), .D(n21696), .Y(n21700)
         );
  OAI22XL U26438 ( .A0(n21705), .A1(n21704), .B0(n22712), .B1(n21703), .Y(
        n21706) );
  AOI21XL U26439 ( .A0(n16663), .A1(n21707), .B0(n21706), .Y(n21723) );
  AOI22XL U26440 ( .A0(conv_1[29]), .A1(n21766), .B0(n21761), .B1(n22722), .Y(
        n21721) );
  AOI22XL U26441 ( .A0(conv_1[419]), .A1(n21763), .B0(conv_1[434]), .B1(n21765), .Y(n21720) );
  AOI22XL U26442 ( .A0(n28324), .A1(n21709), .B0(n21708), .B1(n21736), .Y(
        n21719) );
  OAI22XL U26443 ( .A0(n22721), .A1(n21711), .B0(n33852), .B1(n21710), .Y(
        n21717) );
  INVXL U26444 ( .A(conv_1[404]), .Y(n33273) );
  INVXL U26445 ( .A(conv_1[449]), .Y(n27197) );
  OAI22XL U26446 ( .A0(n33273), .A1(n21731), .B0(n27197), .B1(n17171), .Y(
        n21716) );
  INVXL U26447 ( .A(conv_1[14]), .Y(n27368) );
  OAI22XL U26448 ( .A0(n22720), .A1(n21712), .B0(n27368), .B1(n21730), .Y(
        n21715) );
  OAI22XL U26449 ( .A0(n21713), .A1(n28553), .B0(n28606), .B1(n21556), .Y(
        n21714) );
  NOR4XL U26450 ( .A(n21717), .B(n21716), .C(n21715), .D(n21714), .Y(n21718)
         );
  OAI211XL U26451 ( .A0(n21724), .A1(n16672), .B0(n21723), .C0(n21722), .Y(
        n21789) );
  AOI22XL U26452 ( .A0(conv_1[448]), .A1(n21752), .B0(n21725), .B1(n22767), 
        .Y(n21747) );
  AOI2BB2XL U26453 ( .B0(n21761), .B1(n22771), .A0N(n21726), .A1N(n26285), .Y(
        n21746) );
  AOI22XL U26454 ( .A0(n16665), .A1(n21728), .B0(n18463), .B1(n21727), .Y(
        n21745) );
  INVXL U26455 ( .A(conv_1[223]), .Y(n34681) );
  OAI22XL U26456 ( .A0(n33436), .A1(n21729), .B0(n34681), .B1(n21556), .Y(
        n21743) );
  INVXL U26457 ( .A(conv_1[403]), .Y(n34695) );
  OAI22XL U26458 ( .A0(n34695), .A1(n21731), .B0(n27362), .B1(n21730), .Y(
        n21742) );
  AOI22XL U26459 ( .A0(conv_1[433]), .A1(n21765), .B0(conv_1[238]), .B1(n21764), .Y(n21740) );
  AOI22XL U26460 ( .A0(conv_1[418]), .A1(n21763), .B0(n16663), .B1(n21732), 
        .Y(n21739) );
  AOI22XL U26461 ( .A0(n28366), .A1(n21734), .B0(n21756), .B1(n21733), .Y(
        n21738) );
  AOI22XL U26462 ( .A0(n21736), .A1(n21735), .B0(n22772), .B1(n21753), .Y(
        n21737) );
  NAND4XL U26463 ( .A(n21740), .B(n21739), .C(n21738), .D(n21737), .Y(n21741)
         );
  NOR3XL U26464 ( .A(n21743), .B(n21742), .C(n21741), .Y(n21744) );
  NAND4XL U26465 ( .A(n21747), .B(n21746), .C(n21745), .D(n21744), .Y(n21780)
         );
  AOI22XL U26466 ( .A0(conv_1[402]), .A1(n21749), .B0(conv_1[12]), .B1(n21748), 
        .Y(n21779) );
  AOI22XL U26467 ( .A0(conv_1[447]), .A1(n21752), .B0(n21751), .B1(n21750), 
        .Y(n21778) );
  AOI22XL U26468 ( .A0(n28559), .A1(n21754), .B0(n22735), .B1(n21753), .Y(
        n21777) );
  AOI22XL U26469 ( .A0(n28324), .A1(n21757), .B0(n21756), .B1(n21755), .Y(
        n21758) );
  OAI21XL U26470 ( .A0(n21760), .A1(n21759), .B0(n21758), .Y(n21774) );
  AOI22XL U26471 ( .A0(conv_1[222]), .A1(n21762), .B0(n21761), .B1(n22732), 
        .Y(n21772) );
  AOI22XL U26472 ( .A0(conv_1[237]), .A1(n21764), .B0(conv_1[417]), .B1(n21763), .Y(n21771) );
  AOI22XL U26473 ( .A0(conv_1[27]), .A1(n21766), .B0(conv_1[432]), .B1(n21765), 
        .Y(n21770) );
  AOI22XL U26474 ( .A0(n22847), .A1(n21768), .B0(n16663), .B1(n21767), .Y(
        n21769) );
  NAND4XL U26475 ( .A(n21772), .B(n21771), .C(n21770), .D(n21769), .Y(n21773)
         );
  AOI211XL U26476 ( .A0(n16670), .A1(n21775), .B0(n21774), .C0(n21773), .Y(
        n21776) );
  NAND4XL U26477 ( .A(n21779), .B(n21778), .C(n21777), .D(n21776), .Y(n21783)
         );
  NOR3XL U26478 ( .A(pool[24]), .B(n21780), .C(n21783), .Y(n21788) );
  NAND4XL U26479 ( .A(n21786), .B(n21785), .C(n21784), .D(n21783), .Y(n21787)
         );
  NAND2XL U26480 ( .A(n34815), .B(pool[20]), .Y(n21792) );
  OAI21XL U26481 ( .A0(n21793), .A1(n34815), .B0(n21792), .Y(N29236) );
  INVXL U26482 ( .A(conv_1[269]), .Y(n29233) );
  NAND2XL U26483 ( .A(n30672), .B(conv_1[255]), .Y(n23460) );
  NAND2XL U26484 ( .A(n35272), .B(n23460), .Y(n21794) );
  OAI211XL U26485 ( .A0(n35272), .A1(n23460), .B0(n34422), .C0(n21794), .Y(
        n21796) );
  NOR2X1 U26486 ( .A(n21796), .B(n21798), .Y(n23461) );
  OAI2BB1XL U26487 ( .A0N(n21798), .A1N(n21796), .B0(n21795), .Y(n21797) );
  OAI211XL U26488 ( .A0(n34080), .A1(n21798), .B0(n33067), .C0(n21797), .Y(
        n16207) );
  AOI22XL U26489 ( .A0(n21831), .A1(n24040), .B0(n21801), .B1(n21830), .Y(
        n34920) );
  AOI2BB2XL U26490 ( .B0(n34952), .B1(n34902), .A0N(n24042), .A1N(n21960), .Y(
        n21800) );
  AOI22XL U26491 ( .A0(n16659), .A1(n34907), .B0(n34961), .B1(n34911), .Y(
        n21799) );
  OAI211XL U26492 ( .A0(n21801), .A1(n26409), .B0(n21800), .C0(n21799), .Y(
        n21809) );
  AOI22XL U26493 ( .A0(n21954), .A1(conv_2[390]), .B0(n21991), .B1(n34902), 
        .Y(n21803) );
  AOI22XL U26494 ( .A0(n21887), .A1(conv_2[435]), .B0(conv_2[15]), .B1(n22015), 
        .Y(n21802) );
  OAI211XL U26495 ( .A0(n24006), .A1(n22018), .B0(n21803), .C0(n21802), .Y(
        n21804) );
  AOI211XL U26496 ( .A0(conv_2[420]), .A1(n22021), .B0(n21805), .C0(n21804), 
        .Y(n34917) );
  AOI2BB2XL U26497 ( .B0(n28556), .B1(n34913), .A0N(n34910), .A1N(n34958), .Y(
        n21807) );
  OAI211XL U26498 ( .A0(n34917), .A1(n35135), .B0(n21807), .C0(n21806), .Y(
        n21808) );
  AOI211XL U26499 ( .A0(n23783), .A1(n34920), .B0(n21809), .C0(n21808), .Y(
        n22049) );
  INVXL U26500 ( .A(conv_2[18]), .Y(n23585) );
  AOI22XL U26501 ( .A0(n21990), .A1(conv_2[423]), .B0(n21954), .B1(conv_2[393]), .Y(n21814) );
  INVXL U26502 ( .A(conv_2[408]), .Y(n29425) );
  OAI22XL U26503 ( .A0(n21819), .A1(n22014), .B0(n21810), .B1(n29558), .Y(
        n21811) );
  AOI211XL U26504 ( .A0(n21992), .A1(conv_2[3]), .B0(n21812), .C0(n21811), .Y(
        n21813) );
  OAI211XL U26505 ( .A0(n23585), .A1(n21953), .B0(n21814), .C0(n21813), .Y(
        n25849) );
  AOI22XL U26506 ( .A0(n16667), .A1(n25840), .B0(n35234), .B1(n25839), .Y(
        n21816) );
  NAND2XL U26507 ( .A(n28528), .B(n25834), .Y(n21815) );
  OAI211XL U26508 ( .A0(n19767), .A1(n21817), .B0(n21816), .C0(n21815), .Y(
        n21825) );
  OAI22XL U26509 ( .A0(n25836), .A1(n21960), .B0(n21818), .B1(n21959), .Y(
        n21823) );
  AOI22XL U26510 ( .A0(conv_2[228]), .A1(n21999), .B0(n22011), .B1(n25838), 
        .Y(n21822) );
  INVXL U26511 ( .A(n21819), .Y(n25837) );
  AOI22XL U26512 ( .A0(n16744), .A1(conv_2[213]), .B0(n34952), .B1(n25837), 
        .Y(n21821) );
  NAND4BXL U26513 ( .AN(n21823), .B(n21822), .C(n21821), .D(n21820), .Y(n21824) );
  INVXL U26514 ( .A(pool[52]), .Y(n34870) );
  AOI22XL U26515 ( .A0(n21887), .A1(conv_2[437]), .B0(n21991), .B1(n25855), 
        .Y(n21829) );
  AOI22XL U26516 ( .A0(n16734), .A1(conv_2[407]), .B0(n21954), .B1(conv_2[392]), .Y(n21828) );
  AOI22XL U26517 ( .A0(n21990), .A1(conv_2[422]), .B0(conv_2[17]), .B1(n22015), 
        .Y(n21827) );
  NAND2XL U26518 ( .A(conv_2[2]), .B(n21992), .Y(n21826) );
  NAND4XL U26519 ( .A(n21829), .B(n21828), .C(n21827), .D(n21826), .Y(n25869)
         );
  AOI22XL U26520 ( .A0(n21831), .A1(n25867), .B0(n25857), .B1(n21830), .Y(
        n25852) );
  AOI22XL U26521 ( .A0(n34950), .A1(n25854), .B0(n34952), .B1(n25855), .Y(
        n21832) );
  OAI21XL U26522 ( .A0(n34969), .A1(n25852), .B0(n21832), .Y(n21839) );
  AOI22XL U26523 ( .A0(conv_2[227]), .A1(n21999), .B0(conv_2[212]), .B1(n16744), .Y(n21837) );
  AOI22XL U26524 ( .A0(n16659), .A1(n25860), .B0(n21833), .B1(n25867), .Y(
        n21836) );
  AOI22XL U26525 ( .A0(n34961), .A1(n25850), .B0(n34954), .B1(n25857), .Y(
        n21834) );
  NAND4XL U26526 ( .A(n21837), .B(n21836), .C(n21835), .D(n21834), .Y(n21838)
         );
  AOI22XL U26527 ( .A0(n21990), .A1(conv_2[421]), .B0(n16734), .B1(conv_2[406]), .Y(n21844) );
  AOI22XL U26528 ( .A0(n21954), .A1(conv_2[391]), .B0(n21991), .B1(n25876), 
        .Y(n21843) );
  AOI22XL U26529 ( .A0(n21887), .A1(conv_2[436]), .B0(conv_2[1]), .B1(n21992), 
        .Y(n21842) );
  NAND2XL U26530 ( .A(conv_2[16]), .B(n22015), .Y(n21841) );
  NAND4XL U26531 ( .A(n21844), .B(n21843), .C(n21842), .D(n21841), .Y(n25889)
         );
  AOI22XL U26532 ( .A0(n34952), .A1(n25876), .B0(n22011), .B1(n21845), .Y(
        n21847) );
  NAND2XL U26533 ( .A(conv_2[211]), .B(n16744), .Y(n21846) );
  OAI211XL U26534 ( .A0(n21848), .A1(n18208), .B0(n21847), .C0(n21846), .Y(
        n21855) );
  AOI22XL U26535 ( .A0(conv_2[226]), .A1(n21999), .B0(n34950), .B1(n21849), 
        .Y(n21853) );
  AOI22XL U26536 ( .A0(n34961), .A1(n25881), .B0(n35234), .B1(n25882), .Y(
        n21852) );
  AOI22XL U26537 ( .A0(n16659), .A1(n25880), .B0(n16667), .B1(n25870), .Y(
        n21850) );
  NAND4XL U26538 ( .A(n21853), .B(n21852), .C(n21851), .D(n21850), .Y(n21854)
         );
  AOI222XL U26539 ( .A0(pool[51]), .A1(n34868), .B0(pool[51]), .B1(pool[50]), 
        .C0(n34868), .C1(pool[50]), .Y(n21856) );
  AOI222XL U26540 ( .A0(n34870), .A1(n34869), .B0(n34870), .B1(n21856), .C0(
        n34869), .C1(n21856), .Y(n21857) );
  AOI222XL U26541 ( .A0(pool[53]), .A1(n34873), .B0(pool[53]), .B1(n21857), 
        .C0(n34873), .C1(n21857), .Y(n21975) );
  INVXL U26542 ( .A(pool[54]), .Y(n22189) );
  INVXL U26543 ( .A(conv_2[19]), .Y(n29718) );
  AOI22XL U26544 ( .A0(n21887), .A1(conv_2[439]), .B0(conv_2[4]), .B1(n21992), 
        .Y(n21862) );
  INVXL U26545 ( .A(conv_2[394]), .Y(n29060) );
  OAI22XL U26546 ( .A0(n21944), .A1(n28863), .B0(n16669), .B1(n29060), .Y(
        n21859) );
  AOI211XL U26547 ( .A0(conv_2[424]), .A1(n22021), .B0(n21860), .C0(n21859), 
        .Y(n21861) );
  OAI211XL U26548 ( .A0(n29718), .A1(n21953), .B0(n21862), .C0(n21861), .Y(
        n25946) );
  AOI22XL U26549 ( .A0(n35236), .A1(n21863), .B0(conv_2[229]), .B1(n21999), 
        .Y(n21865) );
  NAND2XL U26550 ( .A(n22011), .B(n25930), .Y(n21864) );
  OAI211XL U26551 ( .A0(n21866), .A1(n21960), .B0(n21865), .C0(n21864), .Y(
        n21872) );
  AOI22XL U26552 ( .A0(n26376), .A1(n25939), .B0(conv_2[214]), .B1(n16744), 
        .Y(n21870) );
  AOI22XL U26553 ( .A0(n16659), .A1(n25931), .B0(n16667), .B1(n25933), .Y(
        n21869) );
  AOI2BB2XL U26554 ( .B0(n35234), .B1(n25937), .A0N(n19767), .A1N(n25943), .Y(
        n21868) );
  NAND4XL U26555 ( .A(n21870), .B(n21869), .C(n21868), .D(n21867), .Y(n21871)
         );
  AOI211XL U26556 ( .A0(n28465), .A1(n25946), .B0(n21872), .C0(n21871), .Y(
        n22188) );
  AOI22XL U26557 ( .A0(n21887), .A1(conv_2[440]), .B0(n21954), .B1(conv_2[395]), .Y(n21876) );
  AOI22XL U26558 ( .A0(n21990), .A1(conv_2[425]), .B0(n21991), .B1(n25897), 
        .Y(n21875) );
  AOI22XL U26559 ( .A0(n16734), .A1(conv_2[410]), .B0(conv_2[20]), .B1(n22015), 
        .Y(n21874) );
  NAND2XL U26560 ( .A(conv_2[5]), .B(n21992), .Y(n21873) );
  NAND4XL U26561 ( .A(n21876), .B(n21875), .C(n21874), .D(n21873), .Y(n25910)
         );
  AOI22XL U26562 ( .A0(conv_2[215]), .A1(n16744), .B0(n22011), .B1(n25898), 
        .Y(n21878) );
  NAND2XL U26563 ( .A(conv_2[230]), .B(n21999), .Y(n21877) );
  OAI211XL U26564 ( .A0(n21879), .A1(n21959), .B0(n21878), .C0(n21877), .Y(
        n21886) );
  AOI2BB2XL U26565 ( .B0(n34952), .B1(n25897), .A0N(n21880), .A1N(n21960), .Y(
        n21884) );
  AOI22XL U26566 ( .A0(n16659), .A1(n25902), .B0(n34961), .B1(n25893), .Y(
        n21883) );
  AOI22XL U26567 ( .A0(n16667), .A1(n25901), .B0(n35234), .B1(n25900), .Y(
        n21882) );
  NAND4XL U26568 ( .A(n21884), .B(n21883), .C(n21882), .D(n21881), .Y(n21885)
         );
  AOI211XL U26569 ( .A0(n28465), .A1(n25910), .B0(n21886), .C0(n21885), .Y(
        n21972) );
  AOI22XL U26570 ( .A0(n21954), .A1(conv_2[396]), .B0(n21991), .B1(n25960), 
        .Y(n21891) );
  AOI22XL U26571 ( .A0(n16734), .A1(conv_2[411]), .B0(n21887), .B1(conv_2[441]), .Y(n21890) );
  AOI22XL U26572 ( .A0(n21990), .A1(conv_2[426]), .B0(conv_2[21]), .B1(n22015), 
        .Y(n21889) );
  NAND2XL U26573 ( .A(conv_2[6]), .B(n21992), .Y(n21888) );
  NAND4XL U26574 ( .A(n21891), .B(n21890), .C(n21889), .D(n21888), .Y(n25966)
         );
  AOI22XL U26575 ( .A0(n16659), .A1(n25952), .B0(n34961), .B1(n25950), .Y(
        n21893) );
  NAND2XL U26576 ( .A(n25956), .B(n24056), .Y(n21892) );
  OAI211XL U26577 ( .A0(n25963), .A1(n28575), .B0(n21893), .C0(n21892), .Y(
        n21900) );
  AOI2BB2XL U26578 ( .B0(conv_2[231]), .B1(n21999), .A0N(n21960), .A1N(n25958), 
        .Y(n21898) );
  AOI22XL U26579 ( .A0(n34952), .A1(n25960), .B0(n22011), .B1(n25949), .Y(
        n21897) );
  AOI22XL U26580 ( .A0(conv_2[216]), .A1(n16744), .B0(n21998), .B1(n21894), 
        .Y(n21896) );
  AOI22XL U26581 ( .A0(n16667), .A1(n25951), .B0(n35234), .B1(n25957), .Y(
        n21895) );
  NAND4XL U26582 ( .A(n21898), .B(n21897), .C(n21896), .D(n21895), .Y(n21899)
         );
  AOI211XL U26583 ( .A0(n28465), .A1(n25966), .B0(n21900), .C0(n21899), .Y(
        n21971) );
  AOI22XL U26584 ( .A0(n21990), .A1(conv_2[427]), .B0(n21887), .B1(conv_2[442]), .Y(n21904) );
  AOI22XL U26585 ( .A0(n21954), .A1(conv_2[397]), .B0(n21991), .B1(n25918), 
        .Y(n21903) );
  AOI22XL U26586 ( .A0(n16734), .A1(conv_2[412]), .B0(conv_2[22]), .B1(n22015), 
        .Y(n21902) );
  NAND2XL U26587 ( .A(conv_2[7]), .B(n21992), .Y(n21901) );
  NAND4XL U26588 ( .A(n21904), .B(n21903), .C(n21902), .D(n21901), .Y(n25929)
         );
  AOI22XL U26589 ( .A0(n34952), .A1(n25918), .B0(n22011), .B1(n25911), .Y(
        n21906) );
  NAND2XL U26590 ( .A(conv_2[232]), .B(n21999), .Y(n21905) );
  OAI211XL U26591 ( .A0(n25915), .A1(n21959), .B0(n21906), .C0(n21905), .Y(
        n21912) );
  AOI22XL U26592 ( .A0(conv_2[217]), .A1(n16744), .B0(n34950), .B1(n25912), 
        .Y(n21910) );
  AOI22XL U26593 ( .A0(n16659), .A1(n25919), .B0(n16667), .B1(n25916), .Y(
        n21909) );
  AOI22XL U26594 ( .A0(n34961), .A1(n25921), .B0(n35234), .B1(n25922), .Y(
        n21908) );
  NAND4XL U26595 ( .A(n21910), .B(n21909), .C(n21908), .D(n21907), .Y(n21911)
         );
  AOI211XL U26596 ( .A0(n28465), .A1(n25929), .B0(n21912), .C0(n21911), .Y(
        n21938) );
  AOI22XL U26597 ( .A0(n16659), .A1(n26036), .B0(n34961), .B1(n26035), .Y(
        n21921) );
  AOI22XL U26598 ( .A0(conv_2[220]), .A1(n16744), .B0(n21998), .B1(n21913), 
        .Y(n21920) );
  AOI22XL U26599 ( .A0(n28556), .A1(n26034), .B0(n24056), .B1(n26033), .Y(
        n21919) );
  OAI22XL U26600 ( .A0(n26041), .A1(n28575), .B0(n26040), .B1(n35196), .Y(
        n21917) );
  AOI22XL U26601 ( .A0(n34950), .A1(n21914), .B0(n22011), .B1(n26032), .Y(
        n21915) );
  OAI21XL U26602 ( .A0(n26038), .A1(n22009), .B0(n21915), .Y(n21916) );
  AOI211XL U26603 ( .A0(conv_2[235]), .A1(n21999), .B0(n21917), .C0(n21916), 
        .Y(n21918) );
  NAND4XL U26604 ( .A(n21921), .B(n21920), .C(n21919), .D(n21918), .Y(n22032)
         );
  AOI22XL U26605 ( .A0(n34961), .A1(n26017), .B0(n35234), .B1(n26016), .Y(
        n21924) );
  OAI22XL U26606 ( .A0(n26009), .A1(n21960), .B0(n30437), .B1(n22030), .Y(
        n21922) );
  AOI21XL U26607 ( .A0(n16667), .A1(n26008), .B0(n21922), .Y(n21923) );
  OAI211XL U26608 ( .A0(n26014), .A1(n28479), .B0(n21924), .C0(n21923), .Y(
        n21929) );
  AOI22XL U26609 ( .A0(n21998), .A1(n21925), .B0(n22011), .B1(n26007), .Y(
        n21927) );
  AOI22XL U26610 ( .A0(conv_2[236]), .A1(n21999), .B0(n34952), .B1(n26011), 
        .Y(n21926) );
  NAND4BXL U26611 ( .AN(n21929), .B(n21928), .C(n21927), .D(n21926), .Y(n22031) );
  AOI22XL U26612 ( .A0(conv_2[233]), .A1(n21999), .B0(n22011), .B1(n25969), 
        .Y(n21930) );
  OAI21XL U26613 ( .A0(n21931), .A1(n21960), .B0(n21930), .Y(n21937) );
  AOI22XL U26614 ( .A0(n16667), .A1(n25970), .B0(n35234), .B1(n25972), .Y(
        n21935) );
  AOI2BB2XL U26615 ( .B0(n34952), .B1(n25976), .A0N(n19767), .A1N(n25974), .Y(
        n21933) );
  AOI22XL U26616 ( .A0(n34961), .A1(n25971), .B0(conv_2[218]), .B1(n16744), 
        .Y(n21932) );
  NAND4XL U26617 ( .A(n21935), .B(n21934), .C(n21933), .D(n21932), .Y(n21936)
         );
  AOI211XL U26618 ( .A0(n35236), .A1(n25977), .B0(n21937), .C0(n21936), .Y(
        n22035) );
  NAND2XL U26619 ( .A(n22035), .B(n21938), .Y(n21939) );
  NOR4BXL U26620 ( .AN(n22188), .B(n22032), .C(n22031), .D(n21939), .Y(n21970)
         );
  AOI22XL U26621 ( .A0(n21990), .A1(conv_2[429]), .B0(n21954), .B1(conv_2[399]), .Y(n21943) );
  AOI22XL U26622 ( .A0(n16734), .A1(conv_2[414]), .B0(n21887), .B1(conv_2[444]), .Y(n21942) );
  AOI22XL U26623 ( .A0(conv_2[24]), .A1(n22015), .B0(n21991), .B1(n25992), .Y(
        n21941) );
  NAND2XL U26624 ( .A(conv_2[9]), .B(n21992), .Y(n21940) );
  NAND4XL U26625 ( .A(n21943), .B(n21942), .C(n21941), .D(n21940), .Y(n26002)
         );
  INVXL U26626 ( .A(conv_2[10]), .Y(n28789) );
  AOI22XL U26627 ( .A0(n21990), .A1(conv_2[430]), .B0(n21954), .B1(conv_2[400]), .Y(n21948) );
  INVXL U26628 ( .A(conv_2[25]), .Y(n27919) );
  OAI22XL U26629 ( .A0(n26038), .A1(n22014), .B0(n21944), .B1(n36040), .Y(
        n21945) );
  AOI211XL U26630 ( .A0(conv_2[445]), .A1(n21887), .B0(n21946), .C0(n21945), 
        .Y(n21947) );
  OAI211XL U26631 ( .A0(n28789), .A1(n22018), .B0(n21948), .C0(n21947), .Y(
        n26044) );
  INVXL U26632 ( .A(conv_2[23]), .Y(n33622) );
  OAI22XL U26633 ( .A0(n21944), .A1(n30884), .B0(n33622), .B1(n21953), .Y(
        n21952) );
  AOI22XL U26634 ( .A0(n21990), .A1(conv_2[428]), .B0(n21887), .B1(conv_2[443]), .Y(n21950) );
  AOI22XL U26635 ( .A0(n21954), .A1(conv_2[398]), .B0(n21991), .B1(n25976), 
        .Y(n21949) );
  NAND2XL U26636 ( .A(n21950), .B(n21949), .Y(n21951) );
  AOI211XL U26637 ( .A0(conv_2[8]), .A1(n21992), .B0(n21952), .C0(n21951), .Y(
        n25981) );
  AOI22XL U26638 ( .A0(n16734), .A1(conv_2[416]), .B0(n21887), .B1(conv_2[446]), .Y(n21956) );
  AOI22XL U26639 ( .A0(n21954), .A1(conv_2[401]), .B0(n21991), .B1(n26011), 
        .Y(n21955) );
  OAI211XL U26640 ( .A0(n27696), .A1(n22018), .B0(n21956), .C0(n21955), .Y(
        n21957) );
  AOI211XL U26641 ( .A0(conv_2[431]), .A1(n22021), .B0(n21958), .C0(n21957), 
        .Y(n26021) );
  NAND3BXL U26642 ( .AN(n26044), .B(n25981), .C(n26021), .Y(n21968) );
  AOI2BB2XL U26643 ( .B0(n35234), .B1(n25994), .A0N(n25998), .A1N(n28479), .Y(
        n21966) );
  AOI22XL U26644 ( .A0(n34952), .A1(n25992), .B0(n24056), .B1(n25993), .Y(
        n21964) );
  OAI22XL U26645 ( .A0(n25997), .A1(n21959), .B0(n25989), .B1(n26473), .Y(
        n21963) );
  OAI22XL U26646 ( .A0(n25988), .A1(n21960), .B0(n29159), .B1(n22008), .Y(
        n21962) );
  OAI22XL U26647 ( .A0(n25999), .A1(n28577), .B0(n30429), .B1(n22030), .Y(
        n21961) );
  NOR4BXL U26648 ( .AN(n21964), .B(n21963), .C(n21962), .D(n21961), .Y(n21965)
         );
  NAND3XL U26649 ( .A(n21967), .B(n21966), .C(n21965), .Y(n22034) );
  AOI221XL U26650 ( .A0(n26002), .A1(n28465), .B0(n21968), .B1(n16700), .C0(
        n22034), .Y(n21969) );
  NAND4XL U26651 ( .A(n21972), .B(n21971), .C(n21970), .D(n21969), .Y(n21973)
         );
  AOI22XL U26652 ( .A0(n22011), .A1(n25813), .B0(n34952), .B1(n25819), .Y(
        n21989) );
  AOI22XL U26653 ( .A0(n35236), .A1(n21983), .B0(n34950), .B1(n21976), .Y(
        n21988) );
  OAI22XL U26654 ( .A0(n25823), .A1(n28577), .B0(n31126), .B1(n22030), .Y(
        n21977) );
  AOI211XL U26655 ( .A0(n21999), .A1(conv_2[239]), .B0(n21978), .C0(n21977), 
        .Y(n21987) );
  AOI22XL U26656 ( .A0(n21990), .A1(conv_2[434]), .B0(n21887), .B1(conv_2[449]), .Y(n21982) );
  AOI22XL U26657 ( .A0(n16734), .A1(conv_2[419]), .B0(n21954), .B1(conv_2[404]), .Y(n21981) );
  AOI22XL U26658 ( .A0(conv_2[29]), .A1(n22015), .B0(n21991), .B1(n25819), .Y(
        n21980) );
  NAND2XL U26659 ( .A(conv_2[14]), .B(n21992), .Y(n21979) );
  NAND4XL U26660 ( .A(n21982), .B(n21981), .C(n21980), .D(n21979), .Y(n25826)
         );
  NOR2BXL U26661 ( .AN(n25815), .B(n21983), .Y(n25816) );
  OAI22XL U26662 ( .A0(n19767), .A1(n25816), .B0(n25822), .B1(n28575), .Y(
        n21985) );
  OAI22XL U26663 ( .A0(n25814), .A1(n18196), .B0(n25821), .B1(n28479), .Y(
        n21984) );
  AOI211XL U26664 ( .A0(n28465), .A1(n25826), .B0(n21985), .C0(n21984), .Y(
        n21986) );
  NAND4XL U26665 ( .A(n21989), .B(n21988), .C(n21987), .D(n21986), .Y(n22045)
         );
  AOI22XL U26666 ( .A0(n21887), .A1(conv_2[447]), .B0(n21954), .B1(conv_2[402]), .Y(n21996) );
  AOI22XL U26667 ( .A0(n21990), .A1(conv_2[432]), .B0(n16734), .B1(conv_2[417]), .Y(n21995) );
  AOI22XL U26668 ( .A0(conv_2[27]), .A1(n22015), .B0(n21991), .B1(n26067), .Y(
        n21994) );
  NAND2XL U26669 ( .A(conv_2[12]), .B(n21992), .Y(n21993) );
  NAND4XL U26670 ( .A(n21996), .B(n21995), .C(n21994), .D(n21993), .Y(n26078)
         );
  AOI22XL U26671 ( .A0(conv_2[237]), .A1(n21999), .B0(n21998), .B1(n21997), 
        .Y(n22000) );
  OAI2BB1XL U26672 ( .A0N(n34952), .A1N(n26067), .B0(n22000), .Y(n22006) );
  AOI22XL U26673 ( .A0(conv_2[222]), .A1(n16744), .B0(n34950), .B1(n26065), 
        .Y(n22004) );
  AOI22XL U26674 ( .A0(n28528), .A1(n26068), .B0(n34961), .B1(n26058), .Y(
        n22003) );
  AOI22XL U26675 ( .A0(n35234), .A1(n26060), .B0(n24056), .B1(n26070), .Y(
        n22002) );
  NAND4XL U26676 ( .A(n22004), .B(n22003), .C(n22002), .D(n22001), .Y(n22005)
         );
  AOI211XL U26677 ( .A0(n22011), .A1(n26064), .B0(n22006), .C0(n22005), .Y(
        n22007) );
  OAI2BB1XL U26678 ( .A0N(n16700), .A1N(n26078), .B0(n22007), .Y(n22038) );
  OAI22XL U26679 ( .A0(n26087), .A1(n22009), .B0(n22008), .B1(n33094), .Y(
        n22010) );
  AOI21XL U26680 ( .A0(n22011), .A1(n26080), .B0(n22010), .Y(n22029) );
  AOI22XL U26681 ( .A0(n34961), .A1(n26090), .B0(n34950), .B1(n22012), .Y(
        n22013) );
  OAI21XL U26682 ( .A0(n26088), .A1(n28479), .B0(n22013), .Y(n22026) );
  INVXL U26683 ( .A(conv_2[13]), .Y(n27928) );
  AOI22XL U26684 ( .A0(n16734), .A1(conv_2[418]), .B0(n21954), .B1(conv_2[403]), .Y(n22017) );
  AOI22XL U26685 ( .A0(n21887), .A1(conv_2[448]), .B0(conv_2[28]), .B1(n22015), 
        .Y(n22016) );
  OAI211XL U26686 ( .A0(n27928), .A1(n22018), .B0(n22017), .C0(n22016), .Y(
        n22019) );
  AOI211XL U26687 ( .A0(conv_2[433]), .A1(n22021), .B0(n22020), .C0(n22019), 
        .Y(n26096) );
  AOI22XL U26688 ( .A0(n28556), .A1(n26091), .B0(n35234), .B1(n26092), .Y(
        n22024) );
  OAI211XL U26689 ( .A0(n26096), .A1(n35135), .B0(n22024), .C0(n22023), .Y(
        n22025) );
  AOI211XL U26690 ( .A0(n35236), .A1(n22027), .B0(n22026), .C0(n22025), .Y(
        n22028) );
  OAI211XL U26691 ( .A0(n33267), .A1(n22030), .B0(n22029), .C0(n22028), .Y(
        n22039) );
  NOR3XL U26692 ( .A(pool[54]), .B(n22038), .C(n22039), .Y(n22044) );
  INVXL U26693 ( .A(n22031), .Y(n22033) );
  NOR4BBXL U26694 ( .AN(n22034), .BN(n22032), .C(n22035), .D(n22033), .Y(
        n22042) );
  AOI2BB2XL U26695 ( .B0(n26021), .B1(n22033), .A0N(n26044), .A1N(n22032), .Y(
        n22041) );
  OAI2BB1XL U26696 ( .A0N(n25981), .A1N(n22035), .B0(pool[54]), .Y(n22036) );
  NOR4BBXL U26697 ( .AN(n22039), .BN(n22038), .C(n22037), .D(n22036), .Y(
        n22040) );
  OAI211XL U26698 ( .A0(n28465), .A1(n22042), .B0(n22041), .C0(n22040), .Y(
        n22043) );
  NAND2XL U26699 ( .A(n34871), .B(pool[50]), .Y(n22048) );
  OAI21XL U26700 ( .A0(n22049), .A1(n34871), .B0(n22048), .Y(N29266) );
  AOI22XL U26701 ( .A0(n34888), .A1(n22051), .B0(n22050), .B1(n34890), .Y(
        N29284) );
  AOI22XL U26702 ( .A0(n34888), .A1(n22053), .B0(n22052), .B1(n34890), .Y(
        N29285) );
  INVXL U26703 ( .A(filter_2[27]), .Y(n22071) );
  INVXL U26704 ( .A(filter_2[21]), .Y(n22082) );
  AOI22XL U26705 ( .A0(n20603), .A1(n22071), .B0(n22082), .B1(n22105), .Y(
        n14811) );
  INVXL U26706 ( .A(filter_2[38]), .Y(n22067) );
  INVXL U26707 ( .A(filter_2[32]), .Y(n22073) );
  AOI22XL U26708 ( .A0(n36100), .A1(n22067), .B0(n22073), .B1(n22105), .Y(
        n14822) );
  INVXL U26709 ( .A(filter_2[14]), .Y(n22085) );
  INVXL U26710 ( .A(filter_2[8]), .Y(n36098) );
  AOI22XL U26711 ( .A0(n36100), .A1(n22085), .B0(n36098), .B1(n22105), .Y(
        n14798) );
  INVXL U26712 ( .A(filter_2[24]), .Y(n22075) );
  INVXL U26713 ( .A(filter_2[18]), .Y(n22103) );
  AOI22XL U26714 ( .A0(n20603), .A1(n22075), .B0(n22103), .B1(n22105), .Y(
        n14808) );
  INVXL U26715 ( .A(filter_2[45]), .Y(n22059) );
  AOI22XL U26716 ( .A0(n20603), .A1(n22054), .B0(n22059), .B1(n22105), .Y(
        n14835) );
  INVXL U26717 ( .A(filter_2[50]), .Y(n22060) );
  AOI22XL U26718 ( .A0(n20603), .A1(n36142), .B0(n22060), .B1(n22105), .Y(
        n14840) );
  INVXL U26719 ( .A(filter_2[46]), .Y(n22058) );
  AOI22XL U26720 ( .A0(n20603), .A1(n22055), .B0(n22058), .B1(n22105), .Y(
        n14836) );
  INVXL U26721 ( .A(filter_2[49]), .Y(n22056) );
  AOI22XL U26722 ( .A0(n20603), .A1(n36139), .B0(n22056), .B1(n22105), .Y(
        n14839) );
  INVXL U26723 ( .A(filter_2[43]), .Y(n22061) );
  AOI22XL U26724 ( .A0(n20603), .A1(n22056), .B0(n22061), .B1(n22105), .Y(
        n14833) );
  INVXL U26725 ( .A(filter_2[48]), .Y(n22057) );
  AOI22XL U26726 ( .A0(n20603), .A1(n36124), .B0(n22057), .B1(n22105), .Y(
        n14838) );
  INVXL U26727 ( .A(filter_2[42]), .Y(n22062) );
  AOI22XL U26728 ( .A0(n20603), .A1(n22057), .B0(n22062), .B1(n22105), .Y(
        n14832) );
  INVXL U26729 ( .A(filter_2[47]), .Y(n22078) );
  INVXL U26730 ( .A(filter_2[41]), .Y(n22063) );
  AOI22XL U26731 ( .A0(n20603), .A1(n22078), .B0(n22063), .B1(n22105), .Y(
        n14831) );
  INVXL U26732 ( .A(filter_2[40]), .Y(n22064) );
  AOI22XL U26733 ( .A0(n20603), .A1(n22058), .B0(n22064), .B1(n22105), .Y(
        n14830) );
  INVXL U26734 ( .A(filter_2[39]), .Y(n22065) );
  AOI22XL U26735 ( .A0(n20603), .A1(n22059), .B0(n22065), .B1(n22105), .Y(
        n14829) );
  INVXL U26736 ( .A(filter_2[44]), .Y(n22068) );
  AOI22XL U26737 ( .A0(n20603), .A1(n22060), .B0(n22068), .B1(n22105), .Y(
        n14834) );
  INVXL U26738 ( .A(filter_2[37]), .Y(n22066) );
  AOI22XL U26739 ( .A0(n36100), .A1(n22061), .B0(n22066), .B1(n22105), .Y(
        n14827) );
  INVXL U26740 ( .A(filter_2[36]), .Y(n22088) );
  AOI22XL U26741 ( .A0(n36100), .A1(n22062), .B0(n22088), .B1(n22105), .Y(
        n14826) );
  INVXL U26742 ( .A(filter_2[35]), .Y(n22069) );
  AOI22XL U26743 ( .A0(n36100), .A1(n22063), .B0(n22069), .B1(n22105), .Y(
        n14825) );
  INVXL U26744 ( .A(filter_2[34]), .Y(n22070) );
  AOI22XL U26745 ( .A0(n36100), .A1(n22064), .B0(n22070), .B1(n22105), .Y(
        n14824) );
  INVXL U26746 ( .A(filter_2[33]), .Y(n22072) );
  AOI22XL U26747 ( .A0(n36100), .A1(n22065), .B0(n22072), .B1(n22105), .Y(
        n14823) );
  INVXL U26748 ( .A(filter_2[19]), .Y(n22080) );
  INVXL U26749 ( .A(filter_2[13]), .Y(n22104) );
  AOI22XL U26750 ( .A0(n20603), .A1(n22080), .B0(n22104), .B1(n22105), .Y(
        n14803) );
  INVXL U26751 ( .A(filter_2[31]), .Y(n22074) );
  AOI22XL U26752 ( .A0(n36100), .A1(n22066), .B0(n22074), .B1(n22105), .Y(
        n14821) );
  AOI22XL U26753 ( .A0(n20603), .A1(n22068), .B0(n22067), .B1(n22105), .Y(
        n14828) );
  INVXL U26754 ( .A(filter_2[29]), .Y(n22076) );
  AOI22XL U26755 ( .A0(n36100), .A1(n22069), .B0(n22076), .B1(n22105), .Y(
        n14819) );
  INVXL U26756 ( .A(filter_2[28]), .Y(n22077) );
  AOI22XL U26757 ( .A0(n36100), .A1(n22070), .B0(n22077), .B1(n22105), .Y(
        n14818) );
  AOI22XL U26758 ( .A0(n36100), .A1(n22072), .B0(n22071), .B1(n22105), .Y(
        n14817) );
  INVXL U26759 ( .A(filter_2[26]), .Y(n22079) );
  AOI22XL U26760 ( .A0(n36100), .A1(n22073), .B0(n22079), .B1(n22105), .Y(
        n14816) );
  INVXL U26761 ( .A(filter_2[25]), .Y(n22081) );
  AOI22XL U26762 ( .A0(n20603), .A1(n22074), .B0(n22081), .B1(n22105), .Y(
        n14815) );
  INVXL U26763 ( .A(filter_2[30]), .Y(n22087) );
  AOI22XL U26764 ( .A0(n20603), .A1(n22087), .B0(n22075), .B1(n22105), .Y(
        n14814) );
  INVXL U26765 ( .A(filter_2[23]), .Y(n22083) );
  AOI22XL U26766 ( .A0(n20603), .A1(n22076), .B0(n22083), .B1(n22105), .Y(
        n14813) );
  INVXL U26767 ( .A(filter_2[22]), .Y(n22084) );
  AOI22XL U26768 ( .A0(n20603), .A1(n22077), .B0(n22084), .B1(n22105), .Y(
        n14812) );
  INVXL U26769 ( .A(filter_2[53]), .Y(n22099) );
  AOI22XL U26770 ( .A0(n20603), .A1(n22099), .B0(n22078), .B1(n22105), .Y(
        n14837) );
  INVXL U26771 ( .A(filter_2[20]), .Y(n22086) );
  AOI22XL U26772 ( .A0(n20603), .A1(n22079), .B0(n22086), .B1(n22105), .Y(
        n14810) );
  AOI22XL U26773 ( .A0(n20603), .A1(n22081), .B0(n22080), .B1(n22105), .Y(
        n14809) );
  INVXL U26774 ( .A(filter_2[15]), .Y(n22101) );
  AOI22XL U26775 ( .A0(n20603), .A1(n22082), .B0(n22101), .B1(n22105), .Y(
        n14805) );
  INVXL U26776 ( .A(filter_2[17]), .Y(n22100) );
  AOI22XL U26777 ( .A0(n20603), .A1(n22083), .B0(n22100), .B1(n22105), .Y(
        n14807) );
  INVXL U26778 ( .A(filter_2[16]), .Y(n22106) );
  AOI22XL U26779 ( .A0(n20603), .A1(n22084), .B0(n22106), .B1(n22105), .Y(
        n14806) );
  AOI22XL U26780 ( .A0(n20603), .A1(n22086), .B0(n22085), .B1(n22105), .Y(
        n14804) );
  AOI22XL U26781 ( .A0(n36100), .A1(n22088), .B0(n22087), .B1(n22105), .Y(
        n14820) );
  ADDFX1 U26782 ( .A(DP_OP_5170J1_126_4278_n33), .B(DP_OP_5170J1_126_4278_n29), 
        .CI(n22089), .CO(n24564), .S(n20353) );
  AOI22XL U26783 ( .A0(affine_2[28]), .A1(n33367), .B0(n16674), .B1(n22090), 
        .Y(n22091) );
  NAND2XL U26784 ( .A(n22091), .B(n33350), .Y(n16533) );
  ADDFX1 U26785 ( .A(DP_OP_5171J1_127_4278_n33), .B(DP_OP_5171J1_127_4278_n29), 
        .CI(n22092), .CO(n24574), .S(n20183) );
  AOI22XL U26786 ( .A0(affine_2[12]), .A1(n33367), .B0(n16674), .B1(n22093), 
        .Y(n22094) );
  NAND2XL U26787 ( .A(n22094), .B(n33368), .Y(n16567) );
  AOI22XL U26788 ( .A0(n34813), .A1(n22096), .B0(n22095), .B1(n34815), .Y(
        N29240) );
  AOI22XL U26789 ( .A0(n34813), .A1(n22098), .B0(n22097), .B1(n34815), .Y(
        N29239) );
  AOI22XL U26790 ( .A0(n36100), .A1(n36151), .B0(n22099), .B1(n22105), .Y(
        n14843) );
  INVXL U26791 ( .A(filter_2[11]), .Y(n36095) );
  AOI22XL U26792 ( .A0(n36100), .A1(n22100), .B0(n36095), .B1(n22105), .Y(
        n14801) );
  INVXL U26793 ( .A(filter_2[12]), .Y(n22102) );
  INVXL U26794 ( .A(filter_2[6]), .Y(n36094) );
  AOI22XL U26795 ( .A0(n36100), .A1(n22102), .B0(n36094), .B1(n22105), .Y(
        n14796) );
  INVXL U26796 ( .A(filter_2[9]), .Y(n36097) );
  AOI22XL U26797 ( .A0(n36100), .A1(n22101), .B0(n36097), .B1(n22105), .Y(
        n14799) );
  AOI22XL U26798 ( .A0(n36100), .A1(n22103), .B0(n22102), .B1(n22105), .Y(
        n14802) );
  INVXL U26799 ( .A(filter_2[7]), .Y(n36099) );
  AOI22XL U26800 ( .A0(n36100), .A1(n22104), .B0(n36099), .B1(n22105), .Y(
        n14797) );
  INVXL U26801 ( .A(filter_2[10]), .Y(n36096) );
  AOI22XL U26802 ( .A0(n36100), .A1(n22106), .B0(n36096), .B1(n22105), .Y(
        n14800) );
  AOI22XL U26803 ( .A0(n35014), .A1(n22108), .B0(n22107), .B1(n35015), .Y(
        N29330) );
  NAND2XL U26804 ( .A(n30607), .B(conv_3[255]), .Y(n30606) );
  INVXL U26805 ( .A(n30606), .Y(n22109) );
  NAND2XL U26806 ( .A(n22109), .B(n29680), .Y(n22110) );
  NAND2XL U26807 ( .A(n30595), .B(conv_3[256]), .Y(n30594) );
  INVXL U26808 ( .A(n22111), .Y(n22112) );
  XOR2XL U26809 ( .A(n28723), .B(n28722), .Y(n22115) );
  NAND2XL U26810 ( .A(conv_3[259]), .B(n22115), .Y(n22114) );
  OAI211XL U26811 ( .A0(conv_3[259]), .A1(n22115), .B0(n35336), .C0(n22114), 
        .Y(n22116) );
  OAI211XL U26812 ( .A0(n35713), .A1(n22117), .B0(n22116), .C0(n34097), .Y(
        n15762) );
  ADDFX1 U26813 ( .A(DP_OP_5166J1_122_9881_n22), .B(DP_OP_5166J1_122_9881_n27), 
        .CI(n22118), .CO(n25068), .S(n20704) );
  AOI22XL U26814 ( .A0(n33563), .A1(n22119), .B0(affine_1[27]), .B1(n25069), 
        .Y(n22120) );
  NAND2XL U26815 ( .A(n22120), .B(n33412), .Y(n16494) );
  INVXL U26816 ( .A(conv_3[194]), .Y(n32212) );
  INVXL U26817 ( .A(n18856), .Y(n22138) );
  INVXL U26818 ( .A(conv_3[184]), .Y(n22137) );
  AOI22XL U26819 ( .A0(n16659), .A1(n22121), .B0(n22847), .B1(n22171), .Y(
        n22127) );
  AOI22XL U26820 ( .A0(n35130), .A1(n22803), .B0(n34827), .B1(n22123), .Y(
        n22125) );
  NAND2XL U26821 ( .A(n28465), .B(n22804), .Y(n22124) );
  NAND2XL U26822 ( .A(conv_3[180]), .B(n29678), .Y(n34702) );
  NAND2XL U26823 ( .A(n34706), .B(n29680), .Y(n22128) );
  AOI211XL U26824 ( .A0(n30536), .A1(n34702), .B0(n34703), .C0(n22129), .Y(
        n27485) );
  INVXL U26825 ( .A(n22129), .Y(n22130) );
  OAI2BB1XL U26826 ( .A0N(conv_3[181]), .A1N(n27485), .B0(n22130), .Y(n23557)
         );
  AOI222XL U26827 ( .A0(n29732), .A1(n29733), .B0(n29732), .B1(conv_3[183]), 
        .C0(n29733), .C1(conv_3[183]), .Y(n22131) );
  INVXL U26828 ( .A(n22131), .Y(n22132) );
  NAND2XL U26829 ( .A(conv_3[184]), .B(n22135), .Y(n22134) );
  OAI211XL U26830 ( .A0(conv_3[184]), .A1(n22135), .B0(n35336), .C0(n22134), 
        .Y(n22136) );
  OAI211XL U26831 ( .A0(n34704), .A1(n22137), .B0(n34097), .C0(n22136), .Y(
        n15767) );
  NAND2XL U26832 ( .A(n27849), .B(n24467), .Y(n22146) );
  NAND2XL U26833 ( .A(n27849), .B(n29677), .Y(n22144) );
  NAND2XL U26834 ( .A(n30842), .B(conv_3[195]), .Y(n30841) );
  INVXL U26835 ( .A(n30841), .Y(n22141) );
  NAND2XL U26836 ( .A(n22141), .B(n29680), .Y(n22142) );
  OAI32XL U26837 ( .A0(n30536), .A1(n27848), .A2(n22141), .B0(n30841), .B1(
        n29680), .Y(n27505) );
  NAND2XL U26838 ( .A(n27505), .B(conv_3[196]), .Y(n27504) );
  NAND2XL U26839 ( .A(n22142), .B(n27504), .Y(n30799) );
  AOI222XL U26840 ( .A0(n30800), .A1(conv_3[197]), .B0(n30800), .B1(n30799), 
        .C0(conv_3[197]), .C1(n30799), .Y(n22143) );
  NAND2XL U26841 ( .A(n22144), .B(n22143), .Y(n29690) );
  OAI21XL U26842 ( .A0(conv_3[198]), .A1(n29689), .B0(n29690), .Y(n22145) );
  NAND2XL U26843 ( .A(n22146), .B(n22145), .Y(n24473) );
  NOR2BXL U26844 ( .AN(n24473), .B(n24474), .Y(n22148) );
  NAND2XL U26845 ( .A(conv_3[199]), .B(n22148), .Y(n22147) );
  OAI211XL U26846 ( .A0(conv_3[199]), .A1(n22148), .B0(n35336), .C0(n22147), 
        .Y(n22149) );
  OAI211XL U26847 ( .A0(n35646), .A1(n22150), .B0(n34097), .C0(n22149), .Y(
        n15766) );
  NAND2XL U26848 ( .A(n23274), .B(n22450), .Y(n22156) );
  NAND2XL U26849 ( .A(n34461), .B(n29677), .Y(n22162) );
  INVXL U26850 ( .A(conv_3[225]), .Y(n25456) );
  NAND2XL U26851 ( .A(n22158), .B(n25454), .Y(n22160) );
  INVXL U26852 ( .A(n25454), .Y(n22159) );
  AOI221XL U26853 ( .A0(n30536), .A1(n22159), .B0(n29680), .B1(n25454), .C0(
        n29136), .Y(n31039) );
  NAND2XL U26854 ( .A(n31039), .B(conv_3[226]), .Y(n31038) );
  NAND2XL U26855 ( .A(n22160), .B(n31038), .Y(n30845) );
  AOI222XL U26856 ( .A0(n30846), .A1(conv_3[227]), .B0(n30846), .B1(n30845), 
        .C0(conv_3[227]), .C1(n30845), .Y(n22161) );
  NAND2XL U26857 ( .A(conv_3[229]), .B(n22166), .Y(n22165) );
  OAI211XL U26858 ( .A0(conv_3[229]), .A1(n22166), .B0(n35336), .C0(n22165), 
        .Y(n22167) );
  OAI211XL U26859 ( .A0(n35676), .A1(n22168), .B0(n34097), .C0(n22167), .Y(
        n15764) );
  INVXL U26860 ( .A(conv_3[154]), .Y(n22187) );
  AOI22XL U26861 ( .A0(n28528), .A1(n22170), .B0(n22847), .B1(n22169), .Y(
        n22176) );
  NAND2XL U26862 ( .A(n28465), .B(n22937), .Y(n22173) );
  NAND2XL U26863 ( .A(n24467), .B(n34579), .Y(n22183) );
  NAND2XL U26864 ( .A(n29677), .B(n34579), .Y(n22181) );
  INVX2 U26865 ( .A(n34579), .Y(n23296) );
  NOR2X1 U26866 ( .A(n27620), .B(n23296), .Y(n34753) );
  NAND2XL U26867 ( .A(n34753), .B(conv_3[150]), .Y(n22177) );
  NAND2XL U26868 ( .A(n22177), .B(n29680), .Y(n22178) );
  NAND2XL U26869 ( .A(n27497), .B(conv_3[151]), .Y(n27496) );
  NAND2XL U26870 ( .A(n22181), .B(n22180), .Y(n29960) );
  NAND2XL U26871 ( .A(conv_3[154]), .B(n22185), .Y(n22184) );
  OAI211XL U26872 ( .A0(conv_3[154]), .A1(n22185), .B0(n35336), .C0(n22184), 
        .Y(n22186) );
  OAI211XL U26873 ( .A0(n34751), .A1(n22187), .B0(n34097), .C0(n22186), .Y(
        n15769) );
  AOI22XL U26874 ( .A0(n34871), .A1(n22189), .B0(n22188), .B1(n34872), .Y(
        N29270) );
  NAND2XL U26875 ( .A(conv_3[469]), .B(n22193), .Y(n22192) );
  OAI211XL U26876 ( .A0(conv_3[469]), .A1(n22193), .B0(n36020), .C0(n22192), 
        .Y(n22194) );
  OAI211XL U26877 ( .A0(n35813), .A1(n22195), .B0(n34097), .C0(n22194), .Y(
        n15748) );
  AOI22XL U26878 ( .A0(n33563), .A1(n22197), .B0(affine_1[17]), .B1(n25243), 
        .Y(n22198) );
  NAND2XL U26879 ( .A(n22198), .B(n33564), .Y(n16484) );
  AOI22XL U26880 ( .A0(n34943), .A1(n22200), .B0(n22199), .B1(n34940), .Y(
        N29302) );
  INVXL U26881 ( .A(conv_1[539]), .Y(n28005) );
  INVXL U26882 ( .A(conv_1[536]), .Y(n22225) );
  AOI22XL U26883 ( .A0(n22362), .A1(n22202), .B0(n21100), .B1(n22201), .Y(
        n22206) );
  AOI22XL U26884 ( .A0(n22369), .A1(n22204), .B0(n22370), .B1(n22203), .Y(
        n22205) );
  AOI22XL U26885 ( .A0(n18463), .A1(n22889), .B0(n26262), .B1(n22399), .Y(
        n22208) );
  AOI22XL U26886 ( .A0(n28366), .A1(n22397), .B0(n26376), .B1(n22843), .Y(
        n22207) );
  OAI211XL U26887 ( .A0(n22209), .A1(n28553), .B0(n22208), .C0(n22207), .Y(
        n22214) );
  AOI222XL U26888 ( .A0(n22212), .A1(n22369), .B0(n22211), .B1(n22370), .C0(
        n22210), .C1(n21100), .Y(n22892) );
  NAND4XL U26889 ( .A(conv_1[525]), .B(n27429), .C(n30672), .D(n34498), .Y(
        n22216) );
  NAND2XL U26890 ( .A(conv_1[525]), .B(n30672), .Y(n33428) );
  AOI211XL U26891 ( .A0(n35272), .A1(n33428), .B0(n33429), .C0(n22215), .Y(
        n30682) );
  NAND2XL U26892 ( .A(conv_1[526]), .B(n30682), .Y(n30681) );
  NAND2XL U26893 ( .A(n22216), .B(n30681), .Y(n22217) );
  NOR2X1 U26894 ( .A(n22218), .B(n22219), .Y(n22220) );
  NOR2BX1 U26895 ( .AN(n26146), .B(conv_1[529]), .Y(n26148) );
  NAND2XL U26896 ( .A(conv_1[530]), .B(n23696), .Y(n22221) );
  NAND2XL U26897 ( .A(n29241), .B(n22222), .Y(n29209) );
  NAND2XL U26898 ( .A(n29236), .B(n29241), .Y(n29208) );
  NAND2XL U26899 ( .A(conv_1[532]), .B(n29208), .Y(n29235) );
  INVXL U26900 ( .A(conv_1[533]), .Y(n29240) );
  AOI21XL U26901 ( .A0(n29215), .A1(conv_1[534]), .B0(n29216), .Y(n29190) );
  NAND2XL U26902 ( .A(n28751), .B(n22223), .Y(n22224) );
  OAI211XL U26903 ( .A0(n33432), .A1(n22225), .B0(n34281), .C0(n22224), .Y(
        n15927) );
  INVXL U26904 ( .A(n35230), .Y(n34982) );
  AOI22XL U26905 ( .A0(n22762), .A1(conv_3[195]), .B0(n16662), .B1(conv_3[210]), .Y(n22229) );
  AOI22XL U26906 ( .A0(n22690), .A1(conv_3[180]), .B0(n16673), .B1(conv_3[225]), .Y(n22228) );
  AOI22XL U26907 ( .A0(n22762), .A1(conv_3[135]), .B0(n22690), .B1(conv_3[120]), .Y(n22231) );
  AOI22XL U26908 ( .A0(n16662), .A1(conv_3[150]), .B0(n18240), .B1(conv_3[165]), .Y(n22230) );
  NAND2XL U26909 ( .A(n22231), .B(n22230), .Y(n35235) );
  AOI22XL U26910 ( .A0(n22362), .A1(n35232), .B0(n21100), .B1(n35235), .Y(
        n22232) );
  NAND2BXL U26911 ( .AN(n22244), .B(n22232), .Y(n25691) );
  AOI22XL U26912 ( .A0(n16662), .A1(conv_3[330]), .B0(n22690), .B1(conv_3[300]), .Y(n22234) );
  AOI222XL U26913 ( .A0(n34951), .A1(n36246), .B0(n22616), .B1(conv_3[420]), 
        .C0(n21011), .C1(conv_3[435]), .Y(n28288) );
  AOI222XL U26914 ( .A0(n22235), .A1(n21688), .B0(n16673), .B1(conv_3[285]), 
        .C0(conv_3[270]), .C1(n25289), .Y(n28285) );
  OAI22XL U26915 ( .A0(n28288), .A1(n25393), .B0(n28285), .B1(n25402), .Y(
        n22239) );
  AOI22XL U26916 ( .A0(n22762), .A1(conv_3[375]), .B0(n16662), .B1(conv_3[390]), .Y(n22237) );
  NAND2XL U26917 ( .A(n22237), .B(n22236), .Y(n28294) );
  OAI2BB2XL U26918 ( .B0(n34982), .B1(n16721), .A0N(n25399), .A1N(n28294), .Y(
        n22238) );
  AOI211XL U26919 ( .A0(n28289), .A1(n28293), .B0(n22239), .C0(n22238), .Y(
        n26159) );
  AOI22XL U26920 ( .A0(n22690), .A1(conv_3[0]), .B0(n18240), .B1(conv_3[45]), 
        .Y(n22241) );
  AOI22XL U26921 ( .A0(n22762), .A1(conv_3[15]), .B0(n16662), .B1(conv_3[30]), 
        .Y(n22240) );
  INVXL U26922 ( .A(conv_3[105]), .Y(n30832) );
  INVXL U26923 ( .A(conv_3[90]), .Y(n30836) );
  OAI2BB2XL U26924 ( .B0(n22612), .B1(n30836), .A0N(n18658), .A1N(conv_3[60]), 
        .Y(n22242) );
  OAI22XL U26925 ( .A0(N18471), .A1(n26159), .B0(n25688), .B1(n34989), .Y(
        n22246) );
  AOI21XL U26926 ( .A0(n28465), .A1(n25691), .B0(n22246), .Y(n22248) );
  NAND2XL U26927 ( .A(n24569), .B(pool[115]), .Y(n22247) );
  OAI21XL U26928 ( .A0(n22248), .A1(n24569), .B0(n22247), .Y(N29331) );
  AOI22XL U26929 ( .A0(n33563), .A1(n22251), .B0(affine_1[8]), .B1(n22250), 
        .Y(n22252) );
  NAND2XL U26930 ( .A(n22252), .B(n33077), .Y(n16505) );
  AOI22XL U26931 ( .A0(n22847), .A1(n22844), .B0(n35181), .B1(n22396), .Y(
        n22255) );
  AOI22XL U26932 ( .A0(n28414), .A1(n22845), .B0(n16745), .B1(n22402), .Y(
        n22254) );
  AOI22XL U26933 ( .A0(n28465), .A1(n23091), .B0(n34827), .B1(n22403), .Y(
        n22253) );
  NAND2XL U26934 ( .A(conv_1[165]), .B(n30672), .Y(n22258) );
  NAND2XL U26935 ( .A(n33497), .B(n27429), .Y(n33063) );
  AOI21XL U26936 ( .A0(n35272), .A1(n22258), .B0(n22257), .Y(n33064) );
  NAND2XL U26937 ( .A(conv_1[166]), .B(n33064), .Y(n33061) );
  NAND2XL U26938 ( .A(n33063), .B(n33061), .Y(n22260) );
  NAND2XL U26939 ( .A(n33403), .B(n22260), .Y(n22259) );
  OAI31XL U26940 ( .A0(n33403), .A1(n22257), .A2(n22260), .B0(n22259), .Y(
        n24492) );
  NAND2XL U26941 ( .A(n22260), .B(n24909), .Y(n22261) );
  OAI2BB1XL U26942 ( .A0N(conv_1[167]), .A1N(n24492), .B0(n22261), .Y(n22433)
         );
  AOI222X1 U26943 ( .A0(conv_1[169]), .A1(n24496), .B0(conv_1[169]), .B1(
        n24497), .C0(n24496), .C1(n24497), .Y(n22262) );
  NAND2XL U26944 ( .A(n27538), .B(n22262), .Y(n35347) );
  INVXL U26945 ( .A(conv_1[179]), .Y(n26671) );
  AOI22XL U26946 ( .A0(n34028), .A1(n22263), .B0(conv_1[171]), .B1(n23915), 
        .Y(n22264) );
  NAND2XL U26947 ( .A(n22264), .B(n34682), .Y(n16292) );
  AOI22X1 U26948 ( .A0(N18471), .A1(n22268), .B0(n22267), .B1(n28467), .Y(
        n22269) );
  INVXL U26949 ( .A(conv_1[322]), .Y(n23326) );
  NAND2XL U26950 ( .A(conv_1[315]), .B(n30672), .Y(n22270) );
  NAND2XL U26951 ( .A(n33860), .B(n27429), .Y(n23981) );
  AOI21XL U26952 ( .A0(n35272), .A1(n22270), .B0(n22269), .Y(n23982) );
  NAND2XL U26953 ( .A(conv_1[316]), .B(n23982), .Y(n22271) );
  NAND2XL U26954 ( .A(n23981), .B(n22271), .Y(n22273) );
  NAND2XL U26955 ( .A(n33403), .B(n22273), .Y(n22272) );
  OAI31XL U26956 ( .A0(n33403), .A1(n22269), .A2(n22273), .B0(n22272), .Y(
        n30494) );
  NAND2XL U26957 ( .A(n22273), .B(n24909), .Y(n22274) );
  OAI31XL U26958 ( .A0(conv_1[320]), .A1(n29383), .A2(conv_1[321]), .B0(n34259), .Y(n23321) );
  AOI21XL U26959 ( .A0(n23326), .A1(n23321), .B0(n29382), .Y(n23315) );
  INVXL U26960 ( .A(conv_1[320]), .Y(n25270) );
  NAND2XL U26961 ( .A(n29385), .B(conv_1[321]), .Y(n23322) );
  AOI21XL U26962 ( .A0(n23316), .A1(conv_1[323]), .B0(n34259), .Y(n23310) );
  INVXL U26963 ( .A(conv_1[329]), .Y(n22930) );
  AOI22XL U26964 ( .A0(n16657), .A1(n22275), .B0(conv_1[325]), .B1(n25268), 
        .Y(n22276) );
  NAND2XL U26965 ( .A(n22276), .B(n16652), .Y(n16138) );
  ADDFXL U26966 ( .A(conv_1[144]), .B(n35339), .CI(n22277), .CO(n26754), .S(
        n22278) );
  AOI22XL U26967 ( .A0(n32611), .A1(n22278), .B0(conv_1[144]), .B1(n35341), 
        .Y(n22279) );
  NAND2XL U26968 ( .A(n22279), .B(n16652), .Y(n16319) );
  INVXL U26969 ( .A(conv_1[173]), .Y(n27543) );
  ADDFXL U26970 ( .A(conv_1[171]), .B(n23923), .CI(n22280), .CO(n27539), .S(
        n22263) );
  OAI21XL U26971 ( .A0(conv_1[172]), .A1(n27539), .B0(n23923), .Y(n27542) );
  AOI31XL U26972 ( .A0(conv_1[172]), .A1(conv_1[173]), .A2(n27539), .B0(n23923), .Y(n23936) );
  AOI22XL U26973 ( .A0(n24378), .A1(n22281), .B0(conv_1[175]), .B1(n23915), 
        .Y(n22282) );
  NAND2XL U26974 ( .A(n22282), .B(n34696), .Y(n16288) );
  NAND2XL U26975 ( .A(conv_1[270]), .B(n30653), .Y(n30652) );
  INVXL U26976 ( .A(n30652), .Y(n22283) );
  NAND2XL U26977 ( .A(n22283), .B(n27429), .Y(n22284) );
  OAI32XL U26978 ( .A0(n22283), .A1(n33994), .A2(n35272), .B0(n27429), .B1(
        n30652), .Y(n30678) );
  NAND2XL U26979 ( .A(conv_1[271]), .B(n30678), .Y(n30677) );
  AND2XL U26980 ( .A(n22284), .B(n30677), .Y(n22285) );
  NAND2XL U26981 ( .A(n24909), .B(n34711), .Y(n22286) );
  AND2XL U26982 ( .A(n22286), .B(n22285), .Y(n30474) );
  NAND2XL U26983 ( .A(n29339), .B(n22287), .Y(n29371) );
  NAND2XL U26984 ( .A(conv_1[275]), .B(n29371), .Y(n29317) );
  INVXL U26985 ( .A(conv_1[276]), .Y(n29321) );
  OAI21XL U26986 ( .A0(conv_1[277]), .A1(n29344), .B0(n29364), .Y(n35421) );
  INVXL U26987 ( .A(conv_1[284]), .Y(n29257) );
  AOI22XL U26988 ( .A0(n16657), .A1(n22288), .B0(conv_1[279]), .B1(n27966), 
        .Y(n22289) );
  NAND2XL U26989 ( .A(n22289), .B(n34281), .Y(n16184) );
  NAND2XL U26990 ( .A(conv_1[225]), .B(n30672), .Y(n22291) );
  INVXL U26991 ( .A(n22292), .Y(n22290) );
  NAND2XL U26992 ( .A(n23951), .B(conv_1[226]), .Y(n23950) );
  NAND2XL U26993 ( .A(n22292), .B(n23950), .Y(n22293) );
  NAND2XL U26994 ( .A(n24909), .B(n22293), .Y(n23890) );
  AOI2BB1XL U26995 ( .A0N(n33403), .A1N(n29136), .B0(n22293), .Y(n22294) );
  INVXL U26996 ( .A(n22294), .Y(n23889) );
  NAND2XL U26997 ( .A(conv_1[227]), .B(n23889), .Y(n22295) );
  AOI222XL U26998 ( .A0(n23364), .A1(conv_1[228]), .B0(n23364), .B1(n23363), 
        .C0(conv_1[228]), .C1(n23363), .Y(n22296) );
  INVXL U26999 ( .A(n22296), .Y(n22297) );
  NOR2X1 U27000 ( .A(n22298), .B(n22297), .Y(n23910) );
  INVXL U27001 ( .A(conv_1[230]), .Y(n22571) );
  INVXL U27002 ( .A(n35404), .Y(n34276) );
  OAI21XL U27003 ( .A0(conv_1[231]), .A1(n29262), .B0(n35404), .Y(n35398) );
  AOI22XL U27004 ( .A0(n34028), .A1(n22300), .B0(conv_1[233]), .B1(n23362), 
        .Y(n22301) );
  NAND2XL U27005 ( .A(n22301), .B(n34682), .Y(n16230) );
  AOI22XL U27006 ( .A0(n32052), .A1(n22303), .B0(conv_1[176]), .B1(n23915), 
        .Y(n22304) );
  NAND2XL U27007 ( .A(n22304), .B(n34696), .Y(n16287) );
  AOI22XL U27008 ( .A0(n34827), .A1(n22936), .B0(n16755), .B1(n22305), .Y(
        n22307) );
  NAND2XL U27009 ( .A(n26470), .B(n22937), .Y(n22306) );
  NOR3XL U27010 ( .A(n33423), .B(n33536), .C(n35272), .Y(n24432) );
  OAI21XL U27011 ( .A0(n33533), .A1(n27429), .B0(n33535), .Y(n24433) );
  AOI2BB1XL U27012 ( .A0N(conv_1[241]), .A1N(n24432), .B0(n24433), .Y(n22309)
         );
  NAND2XL U27013 ( .A(n22309), .B(n33403), .Y(n22308) );
  OAI31XL U27014 ( .A0(n22309), .A1(n33403), .A2(n24021), .B0(n22308), .Y(
        n24385) );
  NAND2XL U27015 ( .A(n22309), .B(n24909), .Y(n22310) );
  OAI2BB1XL U27016 ( .A0N(conv_1[242]), .A1N(n24385), .B0(n22310), .Y(n24271)
         );
  AOI222XL U27017 ( .A0(conv_1[244]), .A1(n24439), .B0(conv_1[244]), .B1(
        n24440), .C0(n24439), .C1(n24440), .Y(n22311) );
  OAI21XL U27018 ( .A0(conv_1[245]), .A1(n23841), .B0(n33663), .Y(n34328) );
  NAND2XL U27019 ( .A(n35414), .B(n22311), .Y(n23842) );
  AOI21XL U27020 ( .A0(conv_1[245]), .A1(n23842), .B0(n33663), .Y(n34329) );
  INVXL U27021 ( .A(conv_1[254]), .Y(n27987) );
  AOI22XL U27022 ( .A0(n16656), .A1(n22312), .B0(conv_1[247]), .B1(n33658), 
        .Y(n22313) );
  NAND2XL U27023 ( .A(n22313), .B(n34682), .Y(n16216) );
  ADDFXL U27024 ( .A(conv_1[305]), .B(n28644), .CI(n22314), .CO(n24153), .S(
        n22315) );
  AOI22XL U27025 ( .A0(n34028), .A1(n22315), .B0(conv_1[305]), .B1(n24151), 
        .Y(n22316) );
  NAND2XL U27026 ( .A(n22316), .B(n34689), .Y(n16158) );
  INVXL U27027 ( .A(conv_1[308]), .Y(n22549) );
  OAI21XL U27028 ( .A0(conv_1[309]), .A1(n28649), .B0(n28644), .Y(n25282) );
  INVXL U27029 ( .A(conv_1[310]), .Y(n25287) );
  AOI21XL U27030 ( .A0(conv_1[309]), .A1(n24163), .B0(n28644), .Y(n25283) );
  AOI22XL U27031 ( .A0(n33982), .A1(n22320), .B0(conv_1[311]), .B1(n24151), 
        .Y(n22321) );
  NAND2XL U27032 ( .A(n22321), .B(n34696), .Y(n16152) );
  AOI22XL U27033 ( .A0(n28407), .A1(pixel[42]), .B0(n22362), .B1(pixel[46]), 
        .Y(n22326) );
  AOI22XL U27034 ( .A0(n28407), .A1(pixel[40]), .B0(n22362), .B1(pixel[44]), 
        .Y(n22323) );
  AOI22XL U27035 ( .A0(n22370), .A1(pixel[8]), .B0(n22369), .B1(pixel[12]), 
        .Y(n22322) );
  OAI2BB1XL U27036 ( .A0N(n22323), .A1N(n22322), .B0(n22368), .Y(n22325) );
  AOI22XL U27037 ( .A0(n22370), .A1(pixel[10]), .B0(n22369), .B1(pixel[14]), 
        .Y(n22324) );
  AOI32XL U27038 ( .A0(n22326), .A1(n22325), .A2(n22324), .B0(n22740), .B1(
        n22325), .Y(n22346) );
  AOI22XL U27039 ( .A0(n28407), .A1(pixel[43]), .B0(n22362), .B1(pixel[47]), 
        .Y(n22331) );
  AOI22XL U27040 ( .A0(n28407), .A1(pixel[41]), .B0(n22362), .B1(pixel[45]), 
        .Y(n22328) );
  AOI22XL U27041 ( .A0(n22370), .A1(pixel[9]), .B0(n22369), .B1(pixel[13]), 
        .Y(n22327) );
  OAI2BB1XL U27042 ( .A0N(n22328), .A1N(n22327), .B0(n22347), .Y(n22330) );
  AOI22XL U27043 ( .A0(n22370), .A1(pixel[11]), .B0(n22369), .B1(pixel[15]), 
        .Y(n22329) );
  AOI32XL U27044 ( .A0(n22331), .A1(n22330), .A2(n22329), .B0(n22716), .B1(
        n22330), .Y(n22345) );
  AOI22XL U27045 ( .A0(n28407), .A1(pixel[35]), .B0(n22362), .B1(pixel[39]), 
        .Y(n22343) );
  AOI22XL U27046 ( .A0(n28407), .A1(pixel[32]), .B0(n22362), .B1(pixel[36]), 
        .Y(n22333) );
  AOI22XL U27047 ( .A0(n22370), .A1(pixel[0]), .B0(n22369), .B1(pixel[4]), .Y(
        n22332) );
  NAND2XL U27048 ( .A(n22333), .B(n22332), .Y(n22340) );
  AOI22XL U27049 ( .A0(n28407), .A1(pixel[34]), .B0(n22362), .B1(pixel[38]), 
        .Y(n22335) );
  AOI22XL U27050 ( .A0(n22370), .A1(pixel[2]), .B0(n22369), .B1(pixel[6]), .Y(
        n22334) );
  AOI21XL U27051 ( .A0(n22335), .A1(n22334), .B0(n22740), .Y(n22339) );
  AOI22XL U27052 ( .A0(n28407), .A1(pixel[33]), .B0(n22362), .B1(pixel[37]), 
        .Y(n22337) );
  AOI22XL U27053 ( .A0(n22370), .A1(pixel[1]), .B0(n22369), .B1(pixel[5]), .Y(
        n22336) );
  AOI21XL U27054 ( .A0(n22337), .A1(n22336), .B0(n18286), .Y(n22338) );
  AOI22XL U27055 ( .A0(n22370), .A1(pixel[3]), .B0(n22369), .B1(pixel[7]), .Y(
        n22341) );
  AOI22XL U27056 ( .A0(n22370), .A1(pixel[27]), .B0(n22369), .B1(pixel[31]), 
        .Y(n22352) );
  AOI22XL U27057 ( .A0(n28407), .A1(pixel[57]), .B0(n22362), .B1(pixel[61]), 
        .Y(n22349) );
  AOI22XL U27058 ( .A0(n22370), .A1(pixel[25]), .B0(n22369), .B1(pixel[29]), 
        .Y(n22348) );
  OAI2BB1XL U27059 ( .A0N(n22349), .A1N(n22348), .B0(n22347), .Y(n22351) );
  AOI22XL U27060 ( .A0(n28407), .A1(pixel[59]), .B0(n22362), .B1(pixel[63]), 
        .Y(n22350) );
  AOI32XL U27061 ( .A0(n22352), .A1(n22351), .A2(n22350), .B0(n22716), .B1(
        n22351), .Y(n22376) );
  AOI22XL U27062 ( .A0(n22370), .A1(pixel[26]), .B0(n22369), .B1(pixel[30]), 
        .Y(n22357) );
  AOI22XL U27063 ( .A0(n28407), .A1(pixel[56]), .B0(n22362), .B1(pixel[60]), 
        .Y(n22354) );
  AOI22XL U27064 ( .A0(n22370), .A1(pixel[24]), .B0(n22369), .B1(pixel[28]), 
        .Y(n22353) );
  OAI2BB1XL U27065 ( .A0N(n22354), .A1N(n22353), .B0(n22368), .Y(n22356) );
  AOI22XL U27066 ( .A0(n28407), .A1(pixel[58]), .B0(n22362), .B1(pixel[62]), 
        .Y(n22355) );
  AOI32XL U27067 ( .A0(n22357), .A1(n22356), .A2(n22355), .B0(n16715), .B1(
        n22356), .Y(n22375) );
  AOI22XL U27068 ( .A0(n28407), .A1(pixel[51]), .B0(n22362), .B1(pixel[55]), 
        .Y(n22373) );
  AOI22XL U27069 ( .A0(n28407), .A1(pixel[48]), .B0(n22362), .B1(pixel[52]), 
        .Y(n22359) );
  AOI22XL U27070 ( .A0(n22370), .A1(pixel[16]), .B0(n22369), .B1(pixel[20]), 
        .Y(n22358) );
  NAND2XL U27071 ( .A(n22359), .B(n22358), .Y(n22367) );
  AOI22XL U27072 ( .A0(n28407), .A1(pixel[50]), .B0(n22362), .B1(pixel[54]), 
        .Y(n22361) );
  AOI22XL U27073 ( .A0(n22370), .A1(pixel[18]), .B0(n22369), .B1(pixel[22]), 
        .Y(n22360) );
  AOI21XL U27074 ( .A0(n22361), .A1(n22360), .B0(n16715), .Y(n22366) );
  AOI22XL U27075 ( .A0(n28407), .A1(pixel[49]), .B0(n22362), .B1(pixel[53]), 
        .Y(n22364) );
  AOI22XL U27076 ( .A0(n22370), .A1(pixel[17]), .B0(n22369), .B1(pixel[21]), 
        .Y(n22363) );
  AOI21XL U27077 ( .A0(n22364), .A1(n22363), .B0(n18286), .Y(n22365) );
  AOI211XL U27078 ( .A0(n22368), .A1(n22367), .B0(n22366), .C0(n22365), .Y(
        n22372) );
  AOI22XL U27079 ( .A0(n22370), .A1(pixel[19]), .B0(n22369), .B1(pixel[23]), 
        .Y(n22371) );
  AOI32XL U27080 ( .A0(n22373), .A1(n22372), .A2(n22371), .B0(n22716), .B1(
        n22372), .Y(n22374) );
  INVXL U27081 ( .A(n27076), .Y(n22379) );
  INVXL U27082 ( .A(conv_1[6]), .Y(n27080) );
  AOI21XL U27083 ( .A0(conv_1[5]), .A1(intadd_2_n1), .B0(n27278), .Y(n27075)
         );
  AOI221XL U27084 ( .A0(n27278), .A1(conv_1[6]), .B0(n22379), .B1(n27080), 
        .C0(n27075), .Y(n27285) );
  OAI2BB1XL U27085 ( .A0N(n27076), .A1N(n27080), .B0(n27278), .Y(n22380) );
  AOI22XL U27086 ( .A0(n34028), .A1(n22381), .B0(conv_1[9]), .B1(n24536), .Y(
        n22382) );
  NAND2XL U27087 ( .A(n22382), .B(n34682), .Y(n16454) );
  AOI22XL U27088 ( .A0(n33778), .A1(n22384), .B0(conv_1[8]), .B1(n24536), .Y(
        n22385) );
  NAND2XL U27089 ( .A(n22385), .B(n16652), .Y(n16455) );
  AOI22XL U27090 ( .A0(n16656), .A1(n22388), .B0(conv_1[273]), .B1(n27966), 
        .Y(n22389) );
  NAND2XL U27091 ( .A(n22389), .B(n32867), .Y(n16190) );
  NAND2XL U27092 ( .A(conv_1[90]), .B(n26695), .Y(n26694) );
  INVXL U27093 ( .A(n26694), .Y(n22390) );
  NAND2XL U27094 ( .A(n22390), .B(n27429), .Y(n22391) );
  OAI32XL U27095 ( .A0(n22390), .A1(n26509), .A2(n35272), .B0(n27429), .B1(
        n26694), .Y(n26699) );
  NAND2XL U27096 ( .A(conv_1[91]), .B(n26699), .Y(n26698) );
  NAND2XL U27097 ( .A(n24909), .B(n34450), .Y(n22393) );
  INVXL U27098 ( .A(conv_1[104]), .Y(n31341) );
  AOI22XL U27099 ( .A0(n34028), .A1(n22394), .B0(conv_1[93]), .B1(n26515), .Y(
        n22395) );
  NAND2XL U27100 ( .A(n22395), .B(n32867), .Y(n16370) );
  AOI22XL U27101 ( .A0(n22847), .A1(n22397), .B0(n35236), .B1(n22396), .Y(
        n22398) );
  OAI2BB1XL U27102 ( .A0N(n28414), .A1N(n22399), .B0(n22398), .Y(n22400) );
  NAND2XL U27103 ( .A(conv_1[75]), .B(n30672), .Y(n22408) );
  NAND2XL U27104 ( .A(n33494), .B(n27429), .Y(n27024) );
  AOI21XL U27105 ( .A0(n35272), .A1(n22408), .B0(n33020), .Y(n27025) );
  NAND2XL U27106 ( .A(conv_1[76]), .B(n27025), .Y(n22409) );
  NAND2XL U27107 ( .A(n27024), .B(n22409), .Y(n22411) );
  NAND2XL U27108 ( .A(n33403), .B(n22411), .Y(n22410) );
  OAI31XL U27109 ( .A0(n33403), .A1(n33020), .A2(n22411), .B0(n22410), .Y(
        n26997) );
  NAND2XL U27110 ( .A(n22411), .B(n24909), .Y(n22412) );
  OAI2BB1XL U27111 ( .A0N(conv_1[77]), .A1N(n26997), .B0(n22412), .Y(n22866)
         );
  AOI22XL U27112 ( .A0(n34028), .A1(n22413), .B0(conv_1[78]), .B1(n24342), .Y(
        n22414) );
  NAND2XL U27113 ( .A(n22414), .B(n32867), .Y(n16385) );
  NAND2XL U27114 ( .A(conv_1[60]), .B(n30672), .Y(n22416) );
  NAND2XL U27115 ( .A(n33488), .B(n27429), .Y(n22417) );
  INVXL U27116 ( .A(n22417), .Y(n22415) );
  AOI211XL U27117 ( .A0(n35272), .A1(n22416), .B0(n31418), .C0(n22415), .Y(
        n27021) );
  NAND2XL U27118 ( .A(conv_1[61]), .B(n27021), .Y(n27020) );
  NAND2XL U27119 ( .A(n24909), .B(n34699), .Y(n22419) );
  AOI22XL U27120 ( .A0(n33982), .A1(n22420), .B0(conv_1[63]), .B1(n33633), .Y(
        n22421) );
  NAND2XL U27121 ( .A(n22421), .B(n32867), .Y(n16400) );
  NAND2XL U27122 ( .A(n30672), .B(conv_1[120]), .Y(n22428) );
  AOI22XL U27123 ( .A0(N18471), .A1(n22422), .B0(n34906), .B1(n23277), .Y(
        n22424) );
  NAND2XL U27124 ( .A(n23785), .B(n23781), .Y(n22423) );
  OAI211XL U27125 ( .A0(n23282), .A1(n34969), .B0(n22424), .C0(n22423), .Y(
        n22425) );
  OR2XL U27126 ( .A(n22428), .B(n28948), .Y(n33491) );
  INVXL U27127 ( .A(conv_1[121]), .Y(n23888) );
  INVXL U27128 ( .A(n28948), .Y(n34493) );
  NAND2XL U27129 ( .A(n35272), .B(n22428), .Y(n22427) );
  OAI211XL U27130 ( .A0(n35272), .A1(n22428), .B0(n34493), .C0(n22427), .Y(
        n23886) );
  OAI21XL U27131 ( .A0(n33403), .A1(n28948), .B0(n30466), .Y(n22430) );
  INVXL U27132 ( .A(n22430), .Y(n30467) );
  INVXL U27133 ( .A(conv_1[122]), .Y(n30472) );
  OAI22XL U27134 ( .A0(n33403), .A1(n30466), .B0(n30467), .B1(n30472), .Y(
        n23647) );
  INVXL U27135 ( .A(conv_1[134]), .Y(n33047) );
  AOI22XL U27136 ( .A0(n33788), .A1(n22431), .B0(conv_1[123]), .B1(n23883), 
        .Y(n22432) );
  NAND2XL U27137 ( .A(n22432), .B(n32867), .Y(n16340) );
  ADDFX1 U27138 ( .A(conv_1[168]), .B(n22434), .CI(n22433), .CO(n24497), .S(
        n22435) );
  AOI22XL U27139 ( .A0(n34028), .A1(n22435), .B0(conv_1[168]), .B1(n23915), 
        .Y(n22436) );
  NAND2XL U27140 ( .A(n22436), .B(n32867), .Y(n16295) );
  AOI22XL U27141 ( .A0(n33778), .A1(n22439), .B0(conv_1[318]), .B1(n25268), 
        .Y(n22440) );
  NAND2XL U27142 ( .A(n22440), .B(n32867), .Y(n16145) );
  INVXL U27143 ( .A(n22443), .Y(n22442) );
  AOI221XL U27144 ( .A0(n22442), .A1(n16656), .B0(n22441), .B1(n34666), .C0(
        n33774), .Y(n22446) );
  AOI31XL U27145 ( .A0(n31735), .A1(n22444), .A2(n22443), .B0(conv_3[451]), 
        .Y(n22445) );
  OAI21XL U27146 ( .A0(n22446), .A1(n22445), .B0(n33550), .Y(n15857) );
  AOI22XL U27147 ( .A0(n23783), .A1(n22450), .B0(n34906), .B1(n22449), .Y(
        n22451) );
  NAND2XL U27148 ( .A(conv_3[45]), .B(n29678), .Y(n23201) );
  INVXL U27149 ( .A(conv_3[59]), .Y(n32184) );
  AOI221XL U27150 ( .A0(n27799), .A1(n32052), .B0(n23201), .B1(n32611), .C0(
        n33818), .Y(n22455) );
  AOI21XL U27151 ( .A0(n34742), .A1(n34507), .B0(conv_3[45]), .Y(n22454) );
  OAI21XL U27152 ( .A0(n22455), .A1(n22454), .B0(n34755), .Y(n15920) );
  INVXL U27153 ( .A(conv_1[411]), .Y(n29291) );
  OAI22XL U27154 ( .A0(n22546), .A1(n23139), .B0(n18321), .B1(n29291), .Y(
        n22457) );
  OAI22XL U27155 ( .A0(n22612), .A1(n29273), .B0(n22717), .B1(n22816), .Y(
        n22456) );
  INVXL U27156 ( .A(conv_1[201]), .Y(n23684) );
  INVXL U27157 ( .A(conv_1[186]), .Y(n35354) );
  OAI22XL U27158 ( .A0(n22546), .A1(n23684), .B0(n22717), .B1(n35354), .Y(
        n22459) );
  OAI22XL U27159 ( .A0(n22612), .A1(n23308), .B0(n24039), .B1(n29267), .Y(
        n22458) );
  OAI22XL U27160 ( .A0(n28500), .A1(n35200), .B0(n28502), .B1(n16672), .Y(
        n22476) );
  AOI222XL U27161 ( .A0(n22460), .A1(n36246), .B0(n22759), .B1(conv_1[426]), 
        .C0(n21011), .C1(conv_1[441]), .Y(n28501) );
  OAI22XL U27162 ( .A0(n19401), .A1(n27349), .B0(n24039), .B1(n27315), .Y(
        n22461) );
  OAI22XL U27163 ( .A0(n28501), .A1(n28349), .B0(n28503), .B1(n35239), .Y(
        n22475) );
  INVXL U27164 ( .A(n25795), .Y(n25771) );
  INVXL U27165 ( .A(conv_1[111]), .Y(n31354) );
  OAI22XL U27166 ( .A0(n22546), .A1(n22871), .B0(n18750), .B1(n31354), .Y(
        n22465) );
  INVXL U27167 ( .A(n28505), .Y(n26586) );
  AOI22XL U27168 ( .A0(n22759), .A1(conv_1[126]), .B0(n16673), .B1(conv_1[171]), .Y(n22467) );
  NAND2XL U27169 ( .A(n22468), .B(n22467), .Y(n28498) );
  AOI22XL U27170 ( .A0(n35236), .A1(n26586), .B0(n16660), .B1(n28498), .Y(
        n22473) );
  AOI22XL U27171 ( .A0(n16716), .A1(conv_1[336]), .B0(n16673), .B1(conv_1[351]), .Y(n22469) );
  NAND2XL U27172 ( .A(n22470), .B(n22469), .Y(n28499) );
  AOI222XL U27173 ( .A0(n22471), .A1(n22765), .B0(n18810), .B1(conv_1[276]), 
        .C0(conv_1[291]), .C1(n16673), .Y(n28504) );
  INVXL U27174 ( .A(n28504), .Y(n26588) );
  AOI22XL U27175 ( .A0(n16665), .A1(n28499), .B0(n28366), .B1(n26588), .Y(
        n22472) );
  OAI211XL U27176 ( .A0(n28511), .A1(n25771), .B0(n22473), .C0(n22472), .Y(
        n22474) );
  NOR3XL U27177 ( .A(n22476), .B(n22475), .C(n22474), .Y(n22789) );
  INVXL U27178 ( .A(conv_1[400]), .Y(n33656) );
  INVXL U27179 ( .A(conv_1[415]), .Y(n29303) );
  OAI22XL U27180 ( .A0(n22612), .A1(n33656), .B0(n24039), .B1(n29303), .Y(
        n22477) );
  AOI211XL U27181 ( .A0(n16666), .A1(conv_1[385]), .B0(n22478), .C0(n22477), 
        .Y(n28454) );
  AOI22XL U27182 ( .A0(n16716), .A1(conv_1[160]), .B0(n22690), .B1(conv_1[130]), .Y(n22479) );
  NAND2XL U27183 ( .A(n22480), .B(n22479), .Y(n28451) );
  INVXL U27184 ( .A(n28451), .Y(n26452) );
  OAI22XL U27185 ( .A0(n28454), .A1(n35200), .B0(n26452), .B1(n35198), .Y(
        n22497) );
  OAI22XL U27186 ( .A0(n22612), .A1(n23009), .B0(n24039), .B1(n28808), .Y(
        n22481) );
  AOI211XL U27187 ( .A0(n22762), .A1(conv_1[325]), .B0(n22482), .C0(n22481), 
        .Y(n28452) );
  INVXL U27188 ( .A(conv_1[220]), .Y(n23295) );
  OAI22XL U27189 ( .A0(n22546), .A1(n35381), .B0(n22717), .B1(n35367), .Y(
        n22483) );
  OAI22XL U27190 ( .A0(n28452), .A1(n28553), .B0(n28456), .B1(n16672), .Y(
        n22496) );
  INVXL U27191 ( .A(conv_1[25]), .Y(n35277) );
  INVXL U27192 ( .A(conv_1[40]), .Y(n35298) );
  INVXL U27193 ( .A(conv_1[55]), .Y(n35318) );
  OAI22XL U27194 ( .A0(n22612), .A1(n35298), .B0(n24039), .B1(n35318), .Y(
        n22485) );
  AOI222XL U27195 ( .A0(n22487), .A1(n21688), .B0(n18810), .B1(conv_1[280]), 
        .C0(conv_1[295]), .C1(n16673), .Y(n28455) );
  INVXL U27196 ( .A(n28455), .Y(n26449) );
  AOI22XL U27197 ( .A0(n28324), .A1(n26449), .B0(n25795), .B1(n28450), .Y(
        n22494) );
  AOI222XL U27198 ( .A0(n22490), .A1(n36246), .B0(n22759), .B1(conv_1[430]), 
        .C0(n22762), .C1(conv_1[445]), .Y(n28453) );
  INVXL U27199 ( .A(n28453), .Y(n24604) );
  INVXL U27200 ( .A(conv_1[70]), .Y(n33640) );
  OAI22XL U27201 ( .A0(n22612), .A1(n26801), .B0(n22717), .B1(n33640), .Y(
        n22491) );
  AOI2BB2XL U27202 ( .B0(n16663), .B1(n24604), .A0N(n18208), .A1N(n28457), .Y(
        n22493) );
  OAI211XL U27203 ( .A0(n28463), .A1(n35239), .B0(n22494), .C0(n22493), .Y(
        n22495) );
  NOR3XL U27204 ( .A(n22497), .B(n22496), .C(n22495), .Y(n22785) );
  INVXL U27205 ( .A(conv_1[274]), .Y(n30771) );
  INVXL U27206 ( .A(conv_1[289]), .Y(n30778) );
  AOI222XL U27207 ( .A0(conv_1[424]), .A1(n22759), .B0(n36246), .B1(n22499), 
        .C0(n25306), .C1(conv_1[439]), .Y(n22500) );
  INVXL U27208 ( .A(n22500), .Y(n25335) );
  AOI22XL U27209 ( .A0(n28324), .A1(n26413), .B0(n16663), .B1(n25335), .Y(
        n22520) );
  AOI22XL U27210 ( .A0(n16662), .A1(conv_1[334]), .B0(n16673), .B1(conv_1[349]), .Y(n22501) );
  NAND2XL U27211 ( .A(n22502), .B(n22501), .Y(n25338) );
  AOI22XL U27212 ( .A0(n16662), .A1(conv_1[394]), .B0(n18658), .B1(conv_1[364]), .Y(n22503) );
  NAND2XL U27213 ( .A(n22504), .B(n22503), .Y(n25339) );
  AOI22XL U27214 ( .A0(n16670), .A1(n25338), .B0(n16664), .B1(n25339), .Y(
        n22519) );
  AOI22XL U27215 ( .A0(n25299), .A1(conv_1[184]), .B0(n16673), .B1(conv_1[229]), .Y(n22505) );
  NAND2XL U27216 ( .A(n22506), .B(n22505), .Y(n26412) );
  AOI22XL U27217 ( .A0(n25299), .A1(conv_1[124]), .B0(n16673), .B1(conv_1[169]), .Y(n22507) );
  NAND2XL U27218 ( .A(n22508), .B(n22507), .Y(n26570) );
  AOI22XL U27219 ( .A0(n22362), .A1(n26412), .B0(n28407), .B1(n26570), .Y(
        n22511) );
  INVXL U27220 ( .A(n26410), .Y(n26411) );
  NAND2XL U27221 ( .A(n16721), .B(n26411), .Y(n22517) );
  NAND2XL U27222 ( .A(n22511), .B(n22517), .Y(n28466) );
  AOI22XL U27223 ( .A0(n22759), .A1(conv_1[64]), .B0(n16673), .B1(conv_1[109]), 
        .Y(n22512) );
  NAND2XL U27224 ( .A(n22513), .B(n22512), .Y(n26569) );
  AOI22XL U27225 ( .A0(n16662), .A1(conv_1[34]), .B0(n16673), .B1(conv_1[49]), 
        .Y(n22515) );
  NAND2XL U27226 ( .A(n22515), .B(n22514), .Y(n25334) );
  AOI22XL U27227 ( .A0(n22362), .A1(n26569), .B0(n28407), .B1(n25334), .Y(
        n22516) );
  NAND2XL U27228 ( .A(n22516), .B(n22517), .Y(n28464) );
  AOI22XL U27229 ( .A0(n35130), .A1(n28466), .B0(n34827), .B1(n28464), .Y(
        n22518) );
  OR2XL U27230 ( .A(n35135), .B(n22517), .Y(n26571) );
  NAND4XL U27231 ( .A(n22520), .B(n22519), .C(n22518), .D(n26571), .Y(n22782)
         );
  INVXL U27232 ( .A(n22782), .Y(n22798) );
  OAI22XL U27233 ( .A0(n22546), .A1(n31112), .B0(n22612), .B1(n34543), .Y(
        n22524) );
  OAI22XL U27234 ( .A0(n22550), .A1(n25064), .B0(n18321), .B1(n35407), .Y(
        n22523) );
  OAI22XL U27235 ( .A0(n28517), .A1(n25771), .B0(n28519), .B1(n16672), .Y(
        n22541) );
  AOI222XL U27236 ( .A0(n22525), .A1(n22765), .B0(n18810), .B1(conv_1[279]), 
        .C0(conv_1[294]), .C1(n16673), .Y(n28518) );
  AOI22XL U27237 ( .A0(n22759), .A1(conv_1[9]), .B0(n16673), .B1(conv_1[54]), 
        .Y(n22527) );
  NAND2XL U27238 ( .A(n22527), .B(n22526), .Y(n28515) );
  OAI2BB2XL U27239 ( .B0(n28518), .B1(n26621), .A0N(n28515), .A1N(n35195), .Y(
        n22540) );
  AOI22XL U27240 ( .A0(n22759), .A1(conv_1[69]), .B0(n16673), .B1(conv_1[114]), 
        .Y(n22529) );
  NAND2XL U27241 ( .A(n22529), .B(n22528), .Y(n28512) );
  INVXL U27242 ( .A(n28512), .Y(n26610) );
  AOI22XL U27243 ( .A0(n16716), .A1(conv_1[399]), .B0(n16673), .B1(conv_1[414]), .Y(n22530) );
  NAND2XL U27244 ( .A(n22531), .B(n22530), .Y(n28513) );
  AOI222XL U27245 ( .A0(n22532), .A1(n36246), .B0(n22759), .B1(conv_1[429]), 
        .C0(n25306), .C1(conv_1[444]), .Y(n28516) );
  INVXL U27246 ( .A(n28516), .Y(n26439) );
  AOI22XL U27247 ( .A0(n16664), .A1(n28513), .B0(n16663), .B1(n26439), .Y(
        n22538) );
  AOI22XL U27248 ( .A0(n22759), .A1(conv_1[129]), .B0(n16673), .B1(conv_1[174]), .Y(n22534) );
  NAND2XL U27249 ( .A(n22534), .B(n22533), .Y(n28514) );
  AOI22XL U27250 ( .A0(n22759), .A1(conv_1[309]), .B0(n16673), .B1(conv_1[354]), .Y(n22535) );
  NAND2XL U27251 ( .A(n22536), .B(n22535), .Y(n28522) );
  AOI22XL U27252 ( .A0(n16660), .A1(n28514), .B0(n16670), .B1(n28522), .Y(
        n22537) );
  OAI211XL U27253 ( .A0(n26610), .A1(n18208), .B0(n22538), .C0(n22537), .Y(
        n22539) );
  NOR3XL U27254 ( .A(n22541), .B(n22540), .C(n22539), .Y(n22784) );
  NAND4XL U27255 ( .A(n22789), .B(n22785), .C(n22798), .D(n22784), .Y(n22705)
         );
  AOI22XL U27256 ( .A0(n16662), .A1(conv_1[158]), .B0(n16673), .B1(conv_1[173]), .Y(n22543) );
  INVXL U27257 ( .A(conv_1[383]), .Y(n35465) );
  INVXL U27258 ( .A(conv_1[368]), .Y(n35457) );
  OAI22XL U27259 ( .A0(n22546), .A1(n35465), .B0(n22717), .B1(n35457), .Y(
        n22545) );
  INVXL U27260 ( .A(conv_1[398]), .Y(n29362) );
  INVXL U27261 ( .A(conv_1[413]), .Y(n27597) );
  OAI22XL U27262 ( .A0(n22612), .A1(n29362), .B0(n18321), .B1(n27597), .Y(
        n22544) );
  OAI22XL U27263 ( .A0(n28440), .A1(n35198), .B0(n28442), .B1(n35200), .Y(
        n22565) );
  INVXL U27264 ( .A(n21011), .Y(n22546) );
  INVXL U27265 ( .A(conv_1[83]), .Y(n24924) );
  INVXL U27266 ( .A(conv_1[98]), .Y(n26788) );
  INVXL U27267 ( .A(conv_1[68]), .Y(n27203) );
  OAI22XL U27268 ( .A0(n22740), .A1(n26788), .B0(n16668), .B1(n27203), .Y(
        n22547) );
  AOI211XL U27269 ( .A0(conv_1[113]), .A1(n16673), .B0(n22548), .C0(n22547), 
        .Y(n28438) );
  INVXL U27270 ( .A(conv_1[338]), .Y(n35436) );
  INVXL U27271 ( .A(conv_1[323]), .Y(n23320) );
  OAI22XL U27272 ( .A0(n19902), .A1(n23320), .B0(n22550), .B1(n22549), .Y(
        n22551) );
  AOI211XL U27273 ( .A0(n16673), .A1(conv_1[353]), .B0(n22552), .C0(n22551), 
        .Y(n28443) );
  OAI22XL U27274 ( .A0(n28438), .A1(n18208), .B0(n28443), .B1(n28553), .Y(
        n22564) );
  INVXL U27275 ( .A(conv_1[53]), .Y(n27321) );
  INVXL U27276 ( .A(conv_1[23]), .Y(n27355) );
  INVXL U27277 ( .A(conv_1[38]), .Y(n27305) );
  OAI22XL U27278 ( .A0(n22546), .A1(n27355), .B0(n22612), .B1(n27305), .Y(
        n22553) );
  AOI211XL U27279 ( .A0(n22759), .A1(conv_1[8]), .B0(n22554), .C0(n22553), .Y(
        n28449) );
  INVXL U27280 ( .A(n28436), .Y(n25346) );
  OAI22XL U27281 ( .A0(n28449), .A1(n35239), .B0(n25346), .B1(n25771), .Y(
        n22563) );
  AOI222XL U27282 ( .A0(n22557), .A1(n22765), .B0(n18810), .B1(conv_1[278]), 
        .C0(conv_1[293]), .C1(n16673), .Y(n28439) );
  AOI22XL U27283 ( .A0(n22759), .A1(conv_1[188]), .B0(n16673), .B1(conv_1[233]), .Y(n22558) );
  NAND2XL U27284 ( .A(n22559), .B(n22558), .Y(n28437) );
  AOI222XL U27285 ( .A0(n22560), .A1(n36246), .B0(n22759), .B1(conv_1[428]), 
        .C0(n16666), .C1(conv_1[443]), .Y(n28441) );
  INVXL U27286 ( .A(n28441), .Y(n25345) );
  AOI22XL U27287 ( .A0(n28559), .A1(n28437), .B0(n16663), .B1(n25345), .Y(
        n22561) );
  OAI21XL U27288 ( .A0(n28439), .A1(n26621), .B0(n22561), .Y(n22562) );
  NOR4XL U27289 ( .A(n22565), .B(n22564), .C(n22563), .D(n22562), .Y(n22780)
         );
  AOI22XL U27290 ( .A0(n16662), .A1(conv_1[335]), .B0(n16673), .B1(conv_1[350]), .Y(n22567) );
  NAND2XL U27291 ( .A(n22567), .B(n22566), .Y(n28485) );
  AOI222XL U27292 ( .A0(n22568), .A1(n36246), .B0(n22690), .B1(conv_1[425]), 
        .C0(n22762), .C1(conv_1[440]), .Y(n28488) );
  INVXL U27293 ( .A(conv_1[50]), .Y(n27325) );
  INVXL U27294 ( .A(conv_1[20]), .Y(n27333) );
  INVXL U27295 ( .A(conv_1[35]), .Y(n27299) );
  OAI22XL U27296 ( .A0(n22546), .A1(n27333), .B0(n22612), .B1(n27299), .Y(
        n22569) );
  AOI211XL U27297 ( .A0(conv_1[5]), .A1(n22759), .B0(n22570), .C0(n22569), .Y(
        n28491) );
  OAI22XL U27298 ( .A0(n28488), .A1(n28349), .B0(n28491), .B1(n35239), .Y(
        n22587) );
  INVXL U27299 ( .A(conv_1[200]), .Y(n23443) );
  INVXL U27300 ( .A(conv_1[185]), .Y(n23592) );
  OAI22XL U27301 ( .A0(n22546), .A1(n23443), .B0(n22717), .B1(n23592), .Y(
        n22572) );
  INVXL U27302 ( .A(n28489), .Y(n26595) );
  AOI22XL U27303 ( .A0(n22616), .A1(conv_1[365]), .B0(n16673), .B1(conv_1[410]), .Y(n22574) );
  NAND2XL U27304 ( .A(n22575), .B(n22574), .Y(n28484) );
  AOI22XL U27305 ( .A0(n28559), .A1(n26595), .B0(n16664), .B1(n28484), .Y(
        n22585) );
  AOI22XL U27306 ( .A0(n16662), .A1(conv_1[95]), .B0(n25299), .B1(conv_1[65]), 
        .Y(n22577) );
  NAND2XL U27307 ( .A(n22577), .B(n22576), .Y(n28486) );
  AOI22XL U27308 ( .A0(n35236), .A1(n28486), .B0(n25795), .B1(n28494), .Y(
        n22584) );
  AOI22XL U27309 ( .A0(n22759), .A1(conv_1[125]), .B0(n16673), .B1(conv_1[170]), .Y(n22580) );
  NAND2XL U27310 ( .A(n22581), .B(n22580), .Y(n28487) );
  AOI222XL U27311 ( .A0(n22582), .A1(n22743), .B0(n18810), .B1(conv_1[275]), 
        .C0(conv_1[290]), .C1(n16673), .Y(n28490) );
  INVXL U27312 ( .A(n28490), .Y(n26594) );
  AOI22XL U27313 ( .A0(n18197), .A1(n28487), .B0(n28324), .B1(n26594), .Y(
        n22583) );
  NAND3XL U27314 ( .A(n22585), .B(n22584), .C(n22583), .Y(n22586) );
  AOI211XL U27315 ( .A0(n16665), .A1(n28485), .B0(n22587), .C0(n22586), .Y(
        n22779) );
  AOI22XL U27316 ( .A0(n22762), .A1(conv_1[326]), .B0(n22759), .B1(conv_1[311]), .Y(n22589) );
  AOI22XL U27317 ( .A0(n16716), .A1(conv_1[341]), .B0(n16673), .B1(conv_1[356]), .Y(n22588) );
  NAND2XL U27318 ( .A(n22589), .B(n22588), .Y(n28527) );
  AOI222XL U27319 ( .A0(n22590), .A1(n36246), .B0(n22759), .B1(conv_1[431]), 
        .C0(n25306), .C1(conv_1[446]), .Y(n28531) );
  INVXL U27320 ( .A(conv_1[221]), .Y(n25441) );
  INVXL U27321 ( .A(conv_1[191]), .Y(n32990) );
  OAI22XL U27322 ( .A0(n22612), .A1(n25441), .B0(n22717), .B1(n32990), .Y(
        n22591) );
  AOI211XL U27323 ( .A0(conv_1[206]), .A1(n25306), .B0(n22592), .C0(n22591), 
        .Y(n28533) );
  OAI22XL U27324 ( .A0(n28531), .A1(n28349), .B0(n28533), .B1(n16672), .Y(
        n22608) );
  AOI22XL U27325 ( .A0(n22762), .A1(conv_1[386]), .B0(n16673), .B1(conv_1[416]), .Y(n22594) );
  AOI22XL U27326 ( .A0(n16716), .A1(conv_1[401]), .B0(n22759), .B1(conv_1[371]), .Y(n22593) );
  NAND2XL U27327 ( .A(n22594), .B(n22593), .Y(n28537) );
  INVXL U27328 ( .A(n28534), .Y(n26444) );
  AOI22XL U27329 ( .A0(n16664), .A1(n28537), .B0(n25795), .B1(n26444), .Y(
        n22606) );
  AOI22XL U27330 ( .A0(n22759), .A1(conv_1[131]), .B0(n16673), .B1(conv_1[176]), .Y(n22597) );
  NAND2XL U27331 ( .A(n22598), .B(n22597), .Y(n28530) );
  AOI222XL U27332 ( .A0(n22599), .A1(n22743), .B0(n18810), .B1(conv_1[281]), 
        .C0(conv_1[296]), .C1(n16673), .Y(n28532) );
  AOI2BB2XL U27333 ( .B0(n16660), .B1(n28530), .A0N(n26621), .A1N(n28532), .Y(
        n22605) );
  AOI22XL U27334 ( .A0(n16716), .A1(conv_1[41]), .B0(n16673), .B1(conv_1[56]), 
        .Y(n22601) );
  AOI22XL U27335 ( .A0(n22762), .A1(conv_1[26]), .B0(n22759), .B1(conv_1[11]), 
        .Y(n22600) );
  NAND2XL U27336 ( .A(n22601), .B(n22600), .Y(n28526) );
  AOI22XL U27337 ( .A0(n16716), .A1(conv_1[101]), .B0(n22690), .B1(conv_1[71]), 
        .Y(n22603) );
  NAND2XL U27338 ( .A(n22603), .B(n22602), .Y(n28529) );
  AOI22XL U27339 ( .A0(n35195), .A1(n28526), .B0(n35236), .B1(n28529), .Y(
        n22604) );
  NAND3XL U27340 ( .A(n22606), .B(n22605), .C(n22604), .Y(n22607) );
  AOI211XL U27341 ( .A0(n16665), .A1(n28527), .B0(n22608), .C0(n22607), .Y(
        n22778) );
  AOI22XL U27342 ( .A0(n16716), .A1(conv_1[157]), .B0(n16673), .B1(conv_1[172]), .Y(n22610) );
  NAND2XL U27343 ( .A(n22610), .B(n22609), .Y(n28475) );
  AOI222XL U27344 ( .A0(n22611), .A1(n36246), .B0(n22690), .B1(conv_1[427]), 
        .C0(n22762), .C1(conv_1[442]), .Y(n28469) );
  INVXL U27345 ( .A(conv_1[202]), .Y(n23450) );
  INVXL U27346 ( .A(conv_1[217]), .Y(n35394) );
  INVXL U27347 ( .A(conv_1[187]), .Y(n23598) );
  OAI22XL U27348 ( .A0(n22612), .A1(n35394), .B0(n22717), .B1(n23598), .Y(
        n22613) );
  OAI22XL U27349 ( .A0(n28469), .A1(n28349), .B0(n28472), .B1(n16672), .Y(
        n22632) );
  AOI22XL U27350 ( .A0(n22616), .A1(conv_1[67]), .B0(n16673), .B1(conv_1[112]), 
        .Y(n22617) );
  NAND2XL U27351 ( .A(n22618), .B(n22617), .Y(n28473) );
  AOI22XL U27352 ( .A0(n22759), .A1(conv_1[367]), .B0(n16673), .B1(conv_1[412]), .Y(n22620) );
  NAND2XL U27353 ( .A(n22620), .B(n22619), .Y(n28474) );
  AOI22XL U27354 ( .A0(n35236), .A1(n28473), .B0(n16664), .B1(n28474), .Y(
        n22630) );
  INVXL U27355 ( .A(conv_1[352]), .Y(n28814) );
  INVXL U27356 ( .A(conv_1[337]), .Y(n23000) );
  OAI22XL U27357 ( .A0(n19902), .A1(n23326), .B0(n22612), .B1(n23000), .Y(
        n22621) );
  AOI211XL U27358 ( .A0(conv_1[307]), .A1(n22759), .B0(n22622), .C0(n22621), 
        .Y(n28480) );
  INVXL U27359 ( .A(n28480), .Y(n24577) );
  AOI222XL U27360 ( .A0(n22623), .A1(n22713), .B0(n18810), .B1(conv_1[277]), 
        .C0(conv_1[292]), .C1(n16673), .Y(n28471) );
  INVXL U27361 ( .A(n28471), .Y(n26579) );
  AOI22XL U27362 ( .A0(n16665), .A1(n24577), .B0(n28366), .B1(n26579), .Y(
        n22629) );
  AOI22XL U27363 ( .A0(n16716), .A1(conv_1[37]), .B0(n25299), .B1(conv_1[7]), 
        .Y(n22625) );
  NAND2XL U27364 ( .A(n22625), .B(n22624), .Y(n28476) );
  INVXL U27365 ( .A(n28470), .Y(n26585) );
  AOI22XL U27366 ( .A0(n35195), .A1(n28476), .B0(n25795), .B1(n26585), .Y(
        n22628) );
  NAND3XL U27367 ( .A(n22630), .B(n22629), .C(n22628), .Y(n22631) );
  AOI211XL U27368 ( .A0(n16660), .A1(n28475), .B0(n22632), .C0(n22631), .Y(
        n22790) );
  NAND4XL U27369 ( .A(n22780), .B(n22779), .C(n22778), .D(n22790), .Y(n22704)
         );
  AOI22XL U27370 ( .A0(n16716), .A1(conv_1[393]), .B0(n22759), .B1(conv_1[363]), .Y(n22634) );
  AOI22XL U27371 ( .A0(n22762), .A1(conv_1[378]), .B0(n16723), .B1(conv_1[408]), .Y(n22633) );
  NAND2XL U27372 ( .A(n22634), .B(n22633), .Y(n25378) );
  AOI222XL U27373 ( .A0(n22635), .A1(n36246), .B0(n22759), .B1(conv_1[423]), 
        .C0(n25306), .C1(conv_1[438]), .Y(n25375) );
  AOI22XL U27374 ( .A0(n16664), .A1(n25378), .B0(n16663), .B1(n24615), .Y(
        n22654) );
  AOI22XL U27375 ( .A0(n22762), .A1(conv_1[318]), .B0(n16662), .B1(conv_1[333]), .Y(n22637) );
  AOI22XL U27376 ( .A0(n22759), .A1(conv_1[303]), .B0(n16673), .B1(conv_1[348]), .Y(n22636) );
  NAND2XL U27377 ( .A(n22637), .B(n22636), .Y(n25380) );
  AOI222XL U27378 ( .A0(n22638), .A1(n22765), .B0(n16673), .B1(conv_1[288]), 
        .C0(conv_1[273]), .C1(n16662), .Y(n25376) );
  INVXL U27379 ( .A(n25376), .Y(n26386) );
  AOI22XL U27380 ( .A0(n16670), .A1(n25380), .B0(n28366), .B1(n26386), .Y(
        n22653) );
  AOI22XL U27381 ( .A0(n22762), .A1(conv_1[198]), .B0(n22616), .B1(conv_1[183]), .Y(n22640) );
  AOI22XL U27382 ( .A0(n16716), .A1(conv_1[213]), .B0(n16673), .B1(conv_1[228]), .Y(n22639) );
  NAND2XL U27383 ( .A(n22640), .B(n22639), .Y(n26385) );
  AOI22XL U27384 ( .A0(n25299), .A1(conv_1[123]), .B0(n16673), .B1(conv_1[168]), .Y(n22642) );
  AOI22XL U27385 ( .A0(n22762), .A1(conv_1[138]), .B0(n16662), .B1(conv_1[153]), .Y(n22641) );
  NAND2XL U27386 ( .A(n22642), .B(n22641), .Y(n26538) );
  AOI22XL U27387 ( .A0(n22362), .A1(n26385), .B0(n28407), .B1(n26538), .Y(
        n22645) );
  NAND2XL U27388 ( .A(n16721), .B(n26384), .Y(n22651) );
  NAND2XL U27389 ( .A(n22645), .B(n22651), .Y(n28426) );
  AOI22XL U27390 ( .A0(n18658), .A1(conv_1[63]), .B0(n16673), .B1(conv_1[108]), 
        .Y(n22647) );
  AOI22XL U27391 ( .A0(n22762), .A1(conv_1[78]), .B0(n16662), .B1(conv_1[93]), 
        .Y(n22646) );
  NAND2XL U27392 ( .A(n22647), .B(n22646), .Y(n26537) );
  AOI22XL U27393 ( .A0(n22762), .A1(conv_1[18]), .B0(n16662), .B1(conv_1[33]), 
        .Y(n22649) );
  AOI22XL U27394 ( .A0(n25299), .A1(conv_1[3]), .B0(n16673), .B1(conv_1[48]), 
        .Y(n22648) );
  NAND2XL U27395 ( .A(n22649), .B(n22648), .Y(n25374) );
  AOI22XL U27396 ( .A0(n22362), .A1(n26537), .B0(n28407), .B1(n25374), .Y(
        n22650) );
  NAND2XL U27397 ( .A(n22650), .B(n22651), .Y(n28425) );
  AOI22XL U27398 ( .A0(n35130), .A1(n28426), .B0(n34827), .B1(n28425), .Y(
        n22652) );
  OR2XL U27399 ( .A(n35241), .B(n22651), .Y(n26539) );
  AOI222XL U27400 ( .A0(n22655), .A1(n22765), .B0(n16673), .B1(conv_1[287]), 
        .C0(conv_1[272]), .C1(n25289), .Y(n26566) );
  AOI22XL U27401 ( .A0(n22762), .A1(conv_1[377]), .B0(n22616), .B1(conv_1[362]), .Y(n22659) );
  AOI22XL U27402 ( .A0(n16716), .A1(conv_1[392]), .B0(n16673), .B1(conv_1[407]), .Y(n22658) );
  NAND2XL U27403 ( .A(n22659), .B(n22658), .Y(n25387) );
  AOI22XL U27404 ( .A0(n28465), .A1(n22673), .B0(n16664), .B1(n25387), .Y(
        n22677) );
  AOI22XL U27405 ( .A0(n16716), .A1(conv_1[332]), .B0(n22690), .B1(conv_1[302]), .Y(n22661) );
  AOI22XL U27406 ( .A0(n22762), .A1(conv_1[317]), .B0(n16673), .B1(conv_1[347]), .Y(n22660) );
  NAND2XL U27407 ( .A(n22661), .B(n22660), .Y(n25384) );
  AOI222XL U27408 ( .A0(n22662), .A1(n36246), .B0(n18658), .B1(conv_1[422]), 
        .C0(n22770), .C1(conv_1[437]), .Y(n26401) );
  AOI22XL U27409 ( .A0(n22690), .A1(conv_1[2]), .B0(n16673), .B1(conv_1[47]), 
        .Y(n22664) );
  AOI22XL U27410 ( .A0(n22762), .A1(conv_1[17]), .B0(n16662), .B1(conv_1[32]), 
        .Y(n22663) );
  NAND2XL U27411 ( .A(n22664), .B(n22663), .Y(n26398) );
  AOI22XL U27412 ( .A0(n22762), .A1(conv_1[77]), .B0(n16662), .B1(conv_1[92]), 
        .Y(n22666) );
  AOI22XL U27413 ( .A0(n25299), .A1(conv_1[62]), .B0(n16673), .B1(conv_1[107]), 
        .Y(n22665) );
  NAND2XL U27414 ( .A(n22666), .B(n22665), .Y(n26399) );
  INVXL U27415 ( .A(n26399), .Y(n26556) );
  AOI211XL U27416 ( .A0(n21100), .A1(n26398), .B0(n22667), .C0(n22673), .Y(
        n28429) );
  AOI22XL U27417 ( .A0(n25299), .A1(conv_1[122]), .B0(n16673), .B1(conv_1[167]), .Y(n22669) );
  AOI22XL U27418 ( .A0(n22762), .A1(conv_1[137]), .B0(n16662), .B1(conv_1[152]), .Y(n22668) );
  NAND2XL U27419 ( .A(n22669), .B(n22668), .Y(n26563) );
  AOI22XL U27420 ( .A0(n16716), .A1(conv_1[212]), .B0(n16673), .B1(conv_1[227]), .Y(n22671) );
  AOI22XL U27421 ( .A0(n22762), .A1(conv_1[197]), .B0(n22690), .B1(conv_1[182]), .Y(n22670) );
  AOI211XL U27422 ( .A0(n28407), .A1(n26563), .B0(n22673), .C0(n22672), .Y(
        n28430) );
  OAI22XL U27423 ( .A0(n28429), .A1(n26575), .B0(n28430), .B1(n34989), .Y(
        n22674) );
  AOI211XL U27424 ( .A0(n16665), .A1(n25384), .B0(n22675), .C0(n22674), .Y(
        n22676) );
  OAI211XL U27425 ( .A0(n26566), .A1(n26621), .B0(n22677), .C0(n22676), .Y(
        n34837) );
  AOI22XL U27426 ( .A0(n16716), .A1(conv_1[211]), .B0(n16673), .B1(conv_1[226]), .Y(n22679) );
  AOI22XL U27427 ( .A0(n22762), .A1(conv_1[196]), .B0(n22616), .B1(conv_1[181]), .Y(n22678) );
  NAND2XL U27428 ( .A(n22679), .B(n22678), .Y(n26395) );
  AOI22XL U27429 ( .A0(n22762), .A1(conv_1[136]), .B0(n16662), .B1(conv_1[151]), .Y(n22681) );
  AOI22XL U27430 ( .A0(n22759), .A1(conv_1[121]), .B0(n22615), .B1(conv_1[166]), .Y(n22680) );
  NAND2XL U27431 ( .A(n22681), .B(n22680), .Y(n26547) );
  AOI22XL U27432 ( .A0(n22362), .A1(n26395), .B0(n21100), .B1(n26547), .Y(
        n22684) );
  NAND2XL U27433 ( .A(n16721), .B(n25400), .Y(n26549) );
  NAND2XL U27434 ( .A(n22684), .B(n26549), .Y(n28432) );
  AOI22XL U27435 ( .A0(n22762), .A1(conv_1[76]), .B0(n16662), .B1(conv_1[91]), 
        .Y(n22686) );
  AOI22XL U27436 ( .A0(n22759), .A1(conv_1[61]), .B0(n22615), .B1(conv_1[106]), 
        .Y(n22685) );
  NAND2XL U27437 ( .A(n22686), .B(n22685), .Y(n26546) );
  AOI22XL U27438 ( .A0(n22762), .A1(conv_1[16]), .B0(n16662), .B1(conv_1[31]), 
        .Y(n22688) );
  AOI22XL U27439 ( .A0(n22759), .A1(conv_1[1]), .B0(n22615), .B1(conv_1[46]), 
        .Y(n22687) );
  NAND2XL U27440 ( .A(n22688), .B(n22687), .Y(n25392) );
  AOI22XL U27441 ( .A0(n22362), .A1(n26546), .B0(n21100), .B1(n25392), .Y(
        n22689) );
  NAND2XL U27442 ( .A(n22689), .B(n26549), .Y(n28431) );
  AOI22XL U27443 ( .A0(n35130), .A1(n28432), .B0(n34827), .B1(n28431), .Y(
        n22700) );
  AOI22XL U27444 ( .A0(n22762), .A1(conv_1[316]), .B0(n16673), .B1(conv_1[346]), .Y(n22692) );
  AOI222XL U27445 ( .A0(n22693), .A1(n36246), .B0(n22616), .B1(conv_1[421]), 
        .C0(n21011), .C1(conv_1[436]), .Y(n25394) );
  OAI22XL U27446 ( .A0(n25396), .A1(n28553), .B0(n25394), .B1(n28349), .Y(
        n22698) );
  AOI22XL U27447 ( .A0(n22759), .A1(conv_1[361]), .B0(n16673), .B1(conv_1[406]), .Y(n22695) );
  AOI22XL U27448 ( .A0(n22762), .A1(conv_1[376]), .B0(n16662), .B1(conv_1[391]), .Y(n22694) );
  NAND2XL U27449 ( .A(n22695), .B(n22694), .Y(n25398) );
  INVXL U27450 ( .A(n25398), .Y(n24624) );
  AOI222XL U27451 ( .A0(n22696), .A1(n21688), .B0(n16673), .B1(conv_1[286]), 
        .C0(conv_1[271]), .C1(n16662), .Y(n26393) );
  OAI22XL U27452 ( .A0(n24624), .A1(n35200), .B0(n26393), .B1(n26621), .Y(
        n22697) );
  AOI222XL U27453 ( .A0(pool[30]), .A1(pool[31]), .B0(pool[30]), .B1(n34836), 
        .C0(pool[31]), .C1(n34836), .Y(n22701) );
  AOI222XL U27454 ( .A0(n34838), .A1(n34837), .B0(n34838), .B1(n22701), .C0(
        n34837), .C1(n22701), .Y(n22702) );
  AOI222XL U27455 ( .A0(n22796), .A1(pool[33]), .B0(n22796), .B1(n22702), .C0(
        pool[33]), .C1(n22702), .Y(n22703) );
  OAI22XL U27456 ( .A0(n19902), .A1(n33122), .B0(n24039), .B1(n33852), .Y(
        n22707) );
  OAI22XL U27457 ( .A0(n22612), .A1(n28606), .B0(n22550), .B1(n32995), .Y(
        n22706) );
  AOI22XL U27458 ( .A0(n18810), .A1(conv_1[404]), .B0(n16673), .B1(conv_1[419]), .Y(n22709) );
  NAND2XL U27459 ( .A(n22709), .B(n22708), .Y(n28411) );
  AOI22XL U27460 ( .A0(n28559), .A1(n26632), .B0(n16664), .B1(n28411), .Y(
        n22729) );
  OAI22XL U27461 ( .A0(n19902), .A1(n26831), .B0(n16668), .B1(n33047), .Y(
        n22710) );
  AOI211XL U27462 ( .A0(n16723), .A1(conv_1[179]), .B0(n22711), .C0(n22710), 
        .Y(n28417) );
  INVXL U27463 ( .A(n28417), .Y(n25312) );
  INVXL U27464 ( .A(conv_1[299]), .Y(n23162) );
  AOI222XL U27465 ( .A0(n23162), .A1(n16673), .B0(n29257), .B1(n18810), .C0(
        n22713), .C1(n22712), .Y(n28413) );
  AOI22XL U27466 ( .A0(n16660), .A1(n25312), .B0(n28366), .B1(n28413), .Y(
        n22728) );
  AOI22XL U27467 ( .A0(n22759), .A1(conv_1[74]), .B0(n16673), .B1(conv_1[119]), 
        .Y(n22714) );
  NAND2XL U27468 ( .A(n22715), .B(n22714), .Y(n28412) );
  OAI22XL U27469 ( .A0(n22740), .A1(n28828), .B0(n22717), .B1(n24814), .Y(
        n22718) );
  AOI211XL U27470 ( .A0(conv_1[329]), .A1(n22347), .B0(n22719), .C0(n22718), 
        .Y(n28416) );
  OAI22XL U27471 ( .A0(n28416), .A1(n28553), .B0(n26633), .B1(n25771), .Y(
        n22726) );
  AOI222XL U27472 ( .A0(n22722), .A1(n36246), .B0(n22690), .B1(conv_1[434]), 
        .C0(n22762), .C1(conv_1[449]), .Y(n28415) );
  AOI22XL U27473 ( .A0(n16716), .A1(conv_1[44]), .B0(n16673), .B1(conv_1[59]), 
        .Y(n22724) );
  AOI22XL U27474 ( .A0(conv_1[29]), .A1(n22347), .B0(n25299), .B1(conv_1[14]), 
        .Y(n22723) );
  NAND2XL U27475 ( .A(n22724), .B(n22723), .Y(n28410) );
  INVXL U27476 ( .A(n28410), .Y(n26634) );
  OAI22XL U27477 ( .A0(n28415), .A1(n28349), .B0(n26634), .B1(n35239), .Y(
        n22725) );
  AOI211XL U27478 ( .A0(n35236), .A1(n28412), .B0(n22726), .C0(n22725), .Y(
        n22727) );
  NAND3XL U27479 ( .A(n22729), .B(n22728), .C(n22727), .Y(n22793) );
  INVXL U27480 ( .A(conv_1[372]), .Y(n34311) );
  INVXL U27481 ( .A(conv_1[387]), .Y(n33093) );
  INVXL U27482 ( .A(conv_1[402]), .Y(n33269) );
  OAI22XL U27483 ( .A0(n19902), .A1(n33093), .B0(n22612), .B1(n33269), .Y(
        n22730) );
  AOI211XL U27484 ( .A0(n16673), .A1(conv_1[417]), .B0(n22731), .C0(n22730), 
        .Y(n28578) );
  INVXL U27485 ( .A(n28578), .Y(n24644) );
  AOI222XL U27486 ( .A0(n22732), .A1(n36246), .B0(n22690), .B1(conv_1[432]), 
        .C0(n22770), .C1(conv_1[447]), .Y(n28580) );
  AOI2BB2XL U27487 ( .B0(n16664), .B1(n24644), .A0N(n28349), .A1N(n28580), .Y(
        n22752) );
  AOI22XL U27488 ( .A0(n22762), .A1(conv_1[327]), .B0(n16673), .B1(conv_1[357]), .Y(n22734) );
  AOI22XL U27489 ( .A0(n16716), .A1(conv_1[342]), .B0(n22690), .B1(conv_1[312]), .Y(n22733) );
  NAND2XL U27490 ( .A(n22734), .B(n22733), .Y(n28572) );
  AOI222XL U27491 ( .A0(n22735), .A1(n21688), .B0(n18810), .B1(conv_1[282]), 
        .C0(conv_1[297]), .C1(n16673), .Y(n28576) );
  INVXL U27492 ( .A(n28576), .Y(n26640) );
  AOI22XL U27493 ( .A0(n16665), .A1(n28572), .B0(n28366), .B1(n26640), .Y(
        n22751) );
  AOI22XL U27494 ( .A0(n16716), .A1(conv_1[162]), .B0(n25299), .B1(conv_1[132]), .Y(n22737) );
  AOI22XL U27495 ( .A0(n22762), .A1(conv_1[147]), .B0(n16673), .B1(conv_1[177]), .Y(n22736) );
  NAND2XL U27496 ( .A(n22737), .B(n22736), .Y(n28573) );
  AOI22XL U27497 ( .A0(n22762), .A1(conv_1[27]), .B0(n16673), .B1(conv_1[57]), 
        .Y(n22739) );
  AOI22XL U27498 ( .A0(n16716), .A1(conv_1[42]), .B0(n22616), .B1(conv_1[12]), 
        .Y(n22738) );
  NAND2XL U27499 ( .A(n22739), .B(n22738), .Y(n28574) );
  INVXL U27500 ( .A(n28574), .Y(n26641) );
  INVXL U27501 ( .A(conv_1[102]), .Y(n31336) );
  INVXL U27502 ( .A(conv_1[72]), .Y(n26310) );
  OAI22XL U27503 ( .A0(n22740), .A1(n31336), .B0(n22550), .B1(n26310), .Y(
        n22742) );
  INVXL U27504 ( .A(conv_1[87]), .Y(n26736) );
  INVXL U27505 ( .A(conv_1[117]), .Y(n29338) );
  OAI22XL U27506 ( .A0(n19902), .A1(n26736), .B0(n24039), .B1(n29338), .Y(
        n22741) );
  OAI22XL U27507 ( .A0(n26641), .A1(n35239), .B0(n28579), .B1(n18208), .Y(
        n22749) );
  INVXL U27508 ( .A(n28570), .Y(n26642) );
  AOI22XL U27509 ( .A0(n22762), .A1(conv_1[207]), .B0(n16673), .B1(conv_1[237]), .Y(n22747) );
  AOI22XL U27510 ( .A0(n16716), .A1(conv_1[222]), .B0(n22616), .B1(conv_1[192]), .Y(n22746) );
  NAND2XL U27511 ( .A(n22747), .B(n22746), .Y(n28583) );
  INVXL U27512 ( .A(n28583), .Y(n25417) );
  OAI22XL U27513 ( .A0(n26642), .A1(n25771), .B0(n25417), .B1(n16672), .Y(
        n22748) );
  AOI211XL U27514 ( .A0(n16660), .A1(n28573), .B0(n22749), .C0(n22748), .Y(
        n22750) );
  NAND3XL U27515 ( .A(n22752), .B(n22751), .C(n22750), .Y(n22786) );
  AOI22XL U27516 ( .A0(n16716), .A1(conv_1[163]), .B0(n16673), .B1(conv_1[178]), .Y(n22754) );
  AOI22XL U27517 ( .A0(n22762), .A1(conv_1[148]), .B0(n22690), .B1(conv_1[133]), .Y(n22753) );
  NAND2XL U27518 ( .A(n22754), .B(n22753), .Y(n28560) );
  INVXL U27519 ( .A(conv_1[208]), .Y(n33116) );
  OAI22XL U27520 ( .A0(n19902), .A1(n33116), .B0(n22612), .B1(n34681), .Y(
        n22756) );
  INVXL U27521 ( .A(conv_1[193]), .Y(n34122) );
  OAI22XL U27522 ( .A0(n22717), .A1(n34122), .B0(n24039), .B1(n33846), .Y(
        n22755) );
  INVXL U27523 ( .A(n28554), .Y(n24641) );
  AOI22XL U27524 ( .A0(n16660), .A1(n28560), .B0(n28559), .B1(n24641), .Y(
        n22777) );
  AOI22XL U27525 ( .A0(n22759), .A1(conv_1[73]), .B0(n16673), .B1(conv_1[118]), 
        .Y(n22758) );
  AOI22XL U27526 ( .A0(n22762), .A1(conv_1[88]), .B0(n16662), .B1(conv_1[103]), 
        .Y(n22757) );
  NAND2XL U27527 ( .A(n22758), .B(n22757), .Y(n28558) );
  AOI22XL U27528 ( .A0(n22762), .A1(conv_1[328]), .B0(n16662), .B1(conv_1[343]), .Y(n22761) );
  AOI22XL U27529 ( .A0(n22759), .A1(conv_1[313]), .B0(n16673), .B1(conv_1[358]), .Y(n22760) );
  NAND2XL U27530 ( .A(n22761), .B(n22760), .Y(n28557) );
  AOI22XL U27531 ( .A0(n35236), .A1(n28558), .B0(n16670), .B1(n28557), .Y(
        n22776) );
  AOI22XL U27532 ( .A0(n22762), .A1(conv_1[388]), .B0(n25299), .B1(conv_1[373]), .Y(n22764) );
  AOI22XL U27533 ( .A0(n16716), .A1(conv_1[403]), .B0(n16673), .B1(conv_1[418]), .Y(n22763) );
  NAND2XL U27534 ( .A(n22764), .B(n22763), .Y(n28555) );
  INVXL U27535 ( .A(conv_1[58]), .Y(n33048) );
  OAI22XL U27536 ( .A0(n22546), .A1(n33436), .B0(n24039), .B1(n33048), .Y(
        n22768) );
  OAI22XL U27537 ( .A0(n28550), .A1(n25771), .B0(n28552), .B1(n35239), .Y(
        n22774) );
  AOI222XL U27538 ( .A0(n22771), .A1(n36246), .B0(n22759), .B1(conv_1[433]), 
        .C0(n22770), .C1(conv_1[448]), .Y(n28549) );
  AOI222XL U27539 ( .A0(n22772), .A1(n22713), .B0(n18810), .B1(conv_1[283]), 
        .C0(conv_1[298]), .C1(n16673), .Y(n28563) );
  OAI22XL U27540 ( .A0(n28549), .A1(n28349), .B0(n28563), .B1(n26621), .Y(
        n22773) );
  AOI211XL U27541 ( .A0(n16664), .A1(n28555), .B0(n22774), .C0(n22773), .Y(
        n22775) );
  NAND3XL U27542 ( .A(n22777), .B(n22776), .C(n22775), .Y(n22781) );
  NOR3XL U27543 ( .A(pool[34]), .B(n22786), .C(n22781), .Y(n22792) );
  NOR4BXL U27544 ( .AN(n22781), .B(n22780), .C(n22779), .D(n22778), .Y(n22788)
         );
  NAND2XL U27545 ( .A(pool[34]), .B(n22782), .Y(n22783) );
  NOR4BXL U27546 ( .AN(n22786), .B(n22785), .C(n22784), .D(n22783), .Y(n22787)
         );
  NAND4BBXL U27547 ( .AN(n22790), .BN(n22789), .C(n22788), .D(n22787), .Y(
        n22791) );
  AOI22XL U27548 ( .A0(n34839), .A1(n22797), .B0(n22796), .B1(n34835), .Y(
        N29249) );
  AOI22XL U27549 ( .A0(n34839), .A1(n22799), .B0(n22798), .B1(n34835), .Y(
        N29250) );
  INVXL U27550 ( .A(n30057), .Y(n22808) );
  OAI32XL U27551 ( .A0(n22808), .A1(n23504), .A2(n35272), .B0(n27429), .B1(
        n30057), .Y(n30132) );
  AOI222XL U27552 ( .A0(n28965), .A1(n28966), .B0(n28965), .B1(conv_1[363]), 
        .C0(n28966), .C1(conv_1[363]), .Y(n22809) );
  INVXL U27553 ( .A(n22809), .Y(n22810) );
  INVXL U27554 ( .A(conv_1[365]), .Y(n22842) );
  AOI2BB1XL U27555 ( .A0N(n35455), .A1N(n22832), .B0(n22833), .Y(n22814) );
  NAND2XL U27556 ( .A(conv_1[366]), .B(n22814), .Y(n22813) );
  OAI211XL U27557 ( .A0(conv_1[366]), .A1(n22814), .B0(n32181), .C0(n22813), 
        .Y(n22815) );
  OAI211XL U27558 ( .A0(n35458), .A1(n22816), .B0(n34544), .C0(n22815), .Y(
        n16097) );
  NAND4XL U27559 ( .A(conv_1[285]), .B(n27429), .C(n30672), .D(n34455), .Y(
        n22822) );
  NAND2XL U27560 ( .A(conv_1[285]), .B(n30672), .Y(n22821) );
  INVXL U27561 ( .A(n22821), .Y(n33516) );
  AOI221XL U27562 ( .A0(n35272), .A1(n22821), .B0(n27429), .B1(n33516), .C0(
        n31871), .Y(n30686) );
  NAND2XL U27563 ( .A(conv_1[286]), .B(n30686), .Y(n30685) );
  AND2XL U27564 ( .A(n22822), .B(n30685), .Y(n22823) );
  NAND2XL U27565 ( .A(n24909), .B(n34455), .Y(n22824) );
  AND2XL U27566 ( .A(n22824), .B(n22823), .Y(n30480) );
  AOI222XL U27567 ( .A0(n30773), .A1(n30774), .B0(n30773), .B1(conv_1[289]), 
        .C0(n30774), .C1(conv_1[289]), .Y(n22825) );
  AND2XL U27568 ( .A(n22827), .B(n22825), .Y(n29310) );
  INVXL U27569 ( .A(conv_1[290]), .Y(n29315) );
  INVXL U27570 ( .A(n22827), .Y(n34319) );
  AOI21XL U27571 ( .A0(conv_1[291]), .A1(n29377), .B0(n34319), .Y(n23169) );
  AOI21XL U27572 ( .A0(conv_1[293]), .A1(n23176), .B0(n34319), .Y(n23181) );
  OAI2BB1XL U27573 ( .A0N(conv_1[295]), .A1N(n23188), .B0(n22827), .Y(n34320)
         );
  NAND4XL U27574 ( .A(conv_1[296]), .B(conv_1[297]), .C(n22827), .D(n34320), 
        .Y(n23164) );
  INVXL U27575 ( .A(conv_1[297]), .Y(n34326) );
  INVXL U27576 ( .A(conv_1[296]), .Y(n34317) );
  INVXL U27577 ( .A(conv_1[293]), .Y(n23180) );
  OR2XL U27578 ( .A(n22827), .B(n22826), .Y(n23175) );
  NAND2XL U27579 ( .A(n23180), .B(n23175), .Y(n23182) );
  OAI21XL U27580 ( .A0(conv_1[295]), .A1(n23187), .B0(n34319), .Y(n34313) );
  NAND2XL U27581 ( .A(n34317), .B(n34313), .Y(n22828) );
  NAND2XL U27582 ( .A(n34319), .B(n22828), .Y(n34321) );
  NAND3XL U27583 ( .A(n34319), .B(n34326), .C(n34321), .Y(n23163) );
  INVXL U27584 ( .A(conv_1[298]), .Y(n23168) );
  AOI22XL U27585 ( .A0(conv_1[298]), .A1(n23164), .B0(n23163), .B1(n23168), 
        .Y(n22830) );
  NAND2XL U27586 ( .A(conv_1[299]), .B(n22830), .Y(n22829) );
  OAI211XL U27587 ( .A0(conv_1[299]), .A1(n22830), .B0(n33822), .C0(n22829), 
        .Y(n22831) );
  OAI211XL U27588 ( .A0(n33442), .A1(n23162), .B0(n34689), .C0(n22831), .Y(
        n16164) );
  INVXL U27589 ( .A(conv_1[367]), .Y(n27578) );
  NAND2XL U27590 ( .A(conv_1[366]), .B(n22832), .Y(n27577) );
  NAND2XL U27591 ( .A(conv_1[368]), .B(n35454), .Y(n23149) );
  AOI21XL U27592 ( .A0(n31363), .A1(n23149), .B0(n23151), .Y(n22835) );
  NAND2XL U27593 ( .A(conv_1[369]), .B(n22835), .Y(n22834) );
  OAI211XL U27594 ( .A0(conv_1[369]), .A1(n22835), .B0(n33778), .C0(n22834), 
        .Y(n22836) );
  OAI211XL U27595 ( .A0(n35458), .A1(n23150), .B0(n16652), .C0(n22836), .Y(
        n16094) );
  NAND2XL U27596 ( .A(conv_1[365]), .B(n22840), .Y(n22839) );
  OAI211XL U27597 ( .A0(conv_1[365]), .A1(n22840), .B0(n30090), .C0(n22839), 
        .Y(n22841) );
  OAI211XL U27598 ( .A0(n35458), .A1(n22842), .B0(n16652), .C0(n22841), .Y(
        n16098) );
  INVXL U27599 ( .A(conv_2[105]), .Y(n22857) );
  NAND2XL U27600 ( .A(n28465), .B(n22850), .Y(n22851) );
  INVX2 U27601 ( .A(n34717), .Y(n34715) );
  NAND2XL U27602 ( .A(conv_2[105]), .B(n22855), .Y(n23574) );
  OAI211XL U27603 ( .A0(conv_2[105]), .A1(n22855), .B0(n30090), .C0(n23574), 
        .Y(n22856) );
  OAI211XL U27604 ( .A0(n35894), .A1(n22857), .B0(n22856), .C0(n34583), .Y(
        n15376) );
  INVXL U27605 ( .A(conv_3[284]), .Y(n32263) );
  INVXL U27606 ( .A(conv_3[274]), .Y(n22865) );
  NAND2XL U27607 ( .A(n24467), .B(n34711), .Y(n22861) );
  NAND2XL U27608 ( .A(conv_3[270]), .B(n29678), .Y(n22858) );
  AOI221XL U27609 ( .A0(n34710), .A1(n29680), .B0(n22858), .B1(n30536), .C0(
        n33994), .Y(n30641) );
  NAND2XL U27610 ( .A(n34710), .B(n29680), .Y(n22859) );
  OAI2BB1XL U27611 ( .A0N(conv_3[271]), .A1N(n30641), .B0(n22859), .Y(n33023)
         );
  AOI222XL U27612 ( .A0(n23492), .A1(n23493), .B0(n23492), .B1(conv_3[273]), 
        .C0(n23493), .C1(conv_3[273]), .Y(n22860) );
  NAND2XL U27613 ( .A(n22861), .B(n22860), .Y(n26327) );
  NOR2BXL U27614 ( .AN(n26327), .B(n26328), .Y(n22863) );
  NAND2XL U27615 ( .A(conv_3[274]), .B(n22863), .Y(n22862) );
  OAI211XL U27616 ( .A0(conv_3[274]), .A1(n22863), .B0(n34028), .C0(n22862), 
        .Y(n22864) );
  OAI211XL U27617 ( .A0(n34709), .A1(n22865), .B0(n34097), .C0(n22864), .Y(
        n15761) );
  INVXL U27618 ( .A(n24931), .Y(n24932) );
  INVXL U27619 ( .A(conv_1[80]), .Y(n24936) );
  INVXL U27620 ( .A(n34053), .Y(n26735) );
  AOI33XL U27621 ( .A0(n34053), .A1(n24932), .A2(n24936), .B0(n24931), .B1(
        conv_1[80]), .B2(n26735), .Y(n22869) );
  OAI2BB1XL U27622 ( .A0N(n22871), .A1N(n22869), .B0(n22868), .Y(n22870) );
  OAI211XL U27623 ( .A0(n34057), .A1(n22871), .B0(n34281), .C0(n22870), .Y(
        n16382) );
  NAND2XL U27624 ( .A(n34450), .B(n29677), .Y(n22875) );
  OR2XL U27625 ( .A(n30833), .B(n30536), .Y(n22873) );
  NAND2XL U27626 ( .A(n27501), .B(conv_3[91]), .Y(n27500) );
  NAND2XL U27627 ( .A(conv_3[94]), .B(n22879), .Y(n22878) );
  OAI211XL U27628 ( .A0(conv_3[94]), .A1(n22879), .B0(n35336), .C0(n22878), 
        .Y(n22880) );
  OAI211XL U27629 ( .A0(n35618), .A1(n22881), .B0(n34097), .C0(n22880), .Y(
        n15773) );
  INVXL U27630 ( .A(conv_2[495]), .Y(n22885) );
  OAI211XL U27631 ( .A0(n22883), .A1(conv_2[495]), .B0(n33982), .C0(n22882), 
        .Y(n22884) );
  OAI211XL U27632 ( .A0(n36091), .A1(n22885), .B0(n34583), .C0(n22884), .Y(
        n15350) );
  NAND2XL U27633 ( .A(n22886), .B(conv_2[465]), .Y(n27859) );
  OAI211XL U27634 ( .A0(n22886), .A1(conv_2[465]), .B0(n33982), .C0(n27859), 
        .Y(n22887) );
  OAI211XL U27635 ( .A0(n34177), .A1(n22888), .B0(n34583), .C0(n22887), .Y(
        n15352) );
  INVXL U27636 ( .A(conv_2[449]), .Y(n27927) );
  INVXL U27637 ( .A(conv_2[435]), .Y(n22895) );
  AOI22XL U27638 ( .A0(n16755), .A1(n23091), .B0(n16670), .B1(n22889), .Y(
        n22891) );
  AOI22XL U27639 ( .A0(n35130), .A1(n23090), .B0(n34827), .B1(n23092), .Y(
        n22890) );
  NAND2XL U27640 ( .A(n22893), .B(conv_2[435]), .Y(n27897) );
  OAI211XL U27641 ( .A0(n22893), .A1(conv_2[435]), .B0(n32052), .C0(n27897), 
        .Y(n22894) );
  OAI211XL U27642 ( .A0(n36070), .A1(n22895), .B0(n34583), .C0(n22894), .Y(
        n15354) );
  INVXL U27643 ( .A(conv_2[139]), .Y(n22905) );
  NAND2XL U27644 ( .A(n28126), .B(n34740), .Y(n22897) );
  NAND2XL U27645 ( .A(conv_2[135]), .B(n28124), .Y(n34425) );
  INVXL U27646 ( .A(conv_2[136]), .Y(n24559) );
  NAND2XL U27647 ( .A(n18913), .B(n34425), .Y(n22898) );
  OAI211XL U27648 ( .A0(n18913), .A1(n34425), .B0(n34740), .C0(n22898), .Y(
        n24557) );
  NAND2XL U27649 ( .A(n28128), .B(n34740), .Y(n34613) );
  INVXL U27650 ( .A(conv_2[137]), .Y(n34620) );
  OR2XL U27651 ( .A(n34613), .B(n34614), .Y(n34615) );
  AOI22XL U27652 ( .A0(n34614), .A1(n34613), .B0(n34620), .B1(n34615), .Y(
        n23037) );
  NAND2XL U27653 ( .A(conv_2[139]), .B(n22903), .Y(n22902) );
  OAI211XL U27654 ( .A0(conv_2[139]), .A1(n22903), .B0(n32052), .C0(n22902), 
        .Y(n22904) );
  OAI211XL U27655 ( .A0(n35902), .A1(n22905), .B0(n34408), .C0(n22904), .Y(
        n15230) );
  NAND2XL U27656 ( .A(n24467), .B(n34717), .Y(n22911) );
  NAND2XL U27657 ( .A(n29677), .B(n34717), .Y(n22909) );
  INVXL U27658 ( .A(n30829), .Y(n22906) );
  NAND2XL U27659 ( .A(n22906), .B(n29680), .Y(n22907) );
  NAND2XL U27660 ( .A(n27520), .B(conv_3[106]), .Y(n27519) );
  AOI222XL U27661 ( .A0(n30794), .A1(conv_3[107]), .B0(n30794), .B1(n30793), 
        .C0(conv_3[107]), .C1(n30793), .Y(n22908) );
  NAND2XL U27662 ( .A(n22909), .B(n22908), .Y(n29651) );
  NAND2XL U27663 ( .A(n22911), .B(n22910), .Y(n31767) );
  NOR2BXL U27664 ( .AN(n31767), .B(n31768), .Y(n22913) );
  NAND2XL U27665 ( .A(conv_3[109]), .B(n22913), .Y(n22912) );
  OAI211XL U27666 ( .A0(conv_3[109]), .A1(n22913), .B0(n35336), .C0(n22912), 
        .Y(n22914) );
  OAI211XL U27667 ( .A0(n34200), .A1(n22915), .B0(n34097), .C0(n22914), .Y(
        n15772) );
  INVXL U27668 ( .A(conv_3[89]), .Y(n32156) );
  INVXL U27669 ( .A(conv_3[79]), .Y(n22925) );
  INVXL U27670 ( .A(conv_3[77]), .Y(n34611) );
  NAND2XL U27671 ( .A(n29680), .B(n34438), .Y(n22916) );
  NAND2XL U27672 ( .A(conv_3[75]), .B(n29678), .Y(n33019) );
  INVXL U27673 ( .A(conv_3[76]), .Y(n24672) );
  NAND2XL U27674 ( .A(n30536), .B(n33019), .Y(n22917) );
  OAI211XL U27675 ( .A0(n30536), .A1(n33019), .B0(n34438), .C0(n22917), .Y(
        n24670) );
  OR2XL U27676 ( .A(n22918), .B(n24668), .Y(n22919) );
  NAND2XL U27677 ( .A(n27619), .B(n22919), .Y(n34606) );
  AOI2BB1XL U27678 ( .A0N(n18997), .A1N(n33020), .B0(n22919), .Y(n34607) );
  AOI21XL U27679 ( .A0(n34611), .A1(n34606), .B0(n34607), .Y(n23729) );
  NAND2XL U27680 ( .A(conv_3[79]), .B(n22923), .Y(n22922) );
  OAI211XL U27681 ( .A0(conv_3[79]), .A1(n22923), .B0(n35336), .C0(n22922), 
        .Y(n22924) );
  OAI211XL U27682 ( .A0(n35610), .A1(n22925), .B0(n34097), .C0(n22924), .Y(
        n15774) );
  NAND4XL U27683 ( .A(conv_1[326]), .B(conv_1[327]), .C(n34258), .D(n29382), 
        .Y(n23328) );
  OR4XL U27684 ( .A(n34258), .B(conv_1[327]), .C(conv_1[326]), .D(n29382), .Y(
        n23327) );
  INVXL U27685 ( .A(conv_1[328]), .Y(n23332) );
  AOI22XL U27686 ( .A0(conv_1[328]), .A1(n23328), .B0(n23327), .B1(n23332), 
        .Y(n22928) );
  NAND2XL U27687 ( .A(conv_1[329]), .B(n22928), .Y(n22927) );
  OAI211XL U27688 ( .A0(conv_1[329]), .A1(n22928), .B0(n27932), .C0(n22927), 
        .Y(n22929) );
  OAI211XL U27689 ( .A0(n33442), .A1(n22930), .B0(n34696), .C0(n22929), .Y(
        n16134) );
  NAND2XL U27690 ( .A(conv_1[105]), .B(n30672), .Y(n34714) );
  NAND2XL U27691 ( .A(n27429), .B(n34717), .Y(n22931) );
  AOI211XL U27692 ( .A0(n35272), .A1(n34714), .B0(n34715), .C0(n22932), .Y(
        n32818) );
  INVXL U27693 ( .A(n22932), .Y(n22933) );
  OAI2BB1XL U27694 ( .A0N(conv_1[106]), .A1N(n32818), .B0(n22933), .Y(n24345)
         );
  INVXL U27695 ( .A(conv_1[119]), .Y(n29261) );
  AOI22XL U27696 ( .A0(n34028), .A1(n22934), .B0(conv_1[107]), .B1(n25090), 
        .Y(n22935) );
  NAND2XL U27697 ( .A(n22935), .B(n33542), .Y(n16356) );
  NAND2XL U27698 ( .A(n28465), .B(n23249), .Y(n22938) );
  NAND2XL U27699 ( .A(conv_1[330]), .B(n30672), .Y(n34521) );
  NAND2XL U27700 ( .A(n27429), .B(n34525), .Y(n22940) );
  AOI211XL U27701 ( .A0(n35272), .A1(n34521), .B0(n34522), .C0(n22941), .Y(
        n23676) );
  INVXL U27702 ( .A(n22941), .Y(n22942) );
  OAI2BB1XL U27703 ( .A0N(conv_1[331]), .A1N(n23676), .B0(n22942), .Y(n22979)
         );
  AOI22XL U27704 ( .A0(n16657), .A1(n22943), .B0(conv_1[332]), .B1(n24242), 
        .Y(n22944) );
  NAND2XL U27705 ( .A(n22944), .B(n33542), .Y(n16131) );
  AOI22XL U27706 ( .A0(n34028), .A1(n22947), .B0(conv_1[304]), .B1(n24151), 
        .Y(n22948) );
  NAND2XL U27707 ( .A(n22948), .B(n35489), .Y(n16159) );
  ADDFXL U27708 ( .A(conv_1[319]), .B(n22950), .CI(n22949), .CO(n29383), .S(
        n22951) );
  AOI22XL U27709 ( .A0(n33788), .A1(n22951), .B0(conv_1[319]), .B1(n25268), 
        .Y(n22952) );
  NAND2XL U27710 ( .A(n22952), .B(n35489), .Y(n16144) );
  ADDFX1 U27711 ( .A(conv_1[79]), .B(n22954), .CI(n22953), .CO(n24931), .S(
        n22955) );
  AOI22XL U27712 ( .A0(n16656), .A1(n22955), .B0(conv_1[79]), .B1(n24342), .Y(
        n22956) );
  NAND2XL U27713 ( .A(n22956), .B(n35489), .Y(n16384) );
  INVXL U27714 ( .A(conv_2[239]), .Y(n33101) );
  NAND3XL U27715 ( .A(n28124), .B(n34461), .C(conv_2[225]), .Y(n22957) );
  INVXL U27716 ( .A(n22957), .Y(n34459) );
  NAND2XL U27717 ( .A(n34459), .B(n28126), .Y(n22958) );
  OAI32XL U27718 ( .A0(n18913), .A1(n34459), .A2(n29136), .B0(n22957), .B1(
        n28126), .Y(n31099) );
  NAND2XL U27719 ( .A(n31099), .B(conv_2[226]), .Y(n31098) );
  NAND2XL U27720 ( .A(n22958), .B(n31098), .Y(n22959) );
  NAND2XL U27721 ( .A(n28128), .B(n22959), .Y(n26934) );
  AOI2BB1XL U27722 ( .A0N(n35853), .A1N(n29136), .B0(n22959), .Y(n22960) );
  INVXL U27723 ( .A(n22960), .Y(n26933) );
  NAND2XL U27724 ( .A(conv_2[227]), .B(n26933), .Y(n22961) );
  XOR2XL U27725 ( .A(n29048), .B(n29047), .Y(n22963) );
  NAND2XL U27726 ( .A(conv_2[228]), .B(n22963), .Y(n22962) );
  OAI211XL U27727 ( .A0(conv_2[228]), .A1(n22963), .B0(n34666), .C0(n22962), 
        .Y(n22964) );
  OAI211XL U27728 ( .A0(n34458), .A1(n22965), .B0(n34105), .C0(n22964), .Y(
        n15260) );
  INVXL U27729 ( .A(conv_2[198]), .Y(n22974) );
  NAND2XL U27730 ( .A(n27849), .B(n28068), .Y(n22970) );
  NAND2XL U27731 ( .A(n34115), .B(conv_2[195]), .Y(n22966) );
  OR2XL U27732 ( .A(n22966), .B(n18913), .Y(n22968) );
  NAND2XL U27733 ( .A(n28126), .B(n22966), .Y(n22967) );
  OAI22XL U27734 ( .A0(n22967), .A1(n27848), .B0(n28126), .B1(n22966), .Y(
        n31095) );
  NAND2XL U27735 ( .A(n31095), .B(conv_2[196]), .Y(n31094) );
  NAND2XL U27736 ( .A(n22968), .B(n31094), .Y(n27415) );
  AOI222XL U27737 ( .A0(n27416), .A1(conv_2[197]), .B0(n27416), .B1(n27415), 
        .C0(conv_2[197]), .C1(n27415), .Y(n22969) );
  NAND2XL U27738 ( .A(n22970), .B(n22969), .Y(n27850) );
  NOR2BXL U27739 ( .AN(n27850), .B(n27851), .Y(n22972) );
  NAND2XL U27740 ( .A(conv_2[198]), .B(n22972), .Y(n22971) );
  OAI211XL U27741 ( .A0(conv_2[198]), .A1(n22972), .B0(n34666), .C0(n22971), 
        .Y(n22973) );
  OAI211XL U27742 ( .A0(n35931), .A1(n22974), .B0(n34105), .C0(n22973), .Y(
        n15262) );
  ADDFX1 U27743 ( .A(conv_1[385]), .B(n35463), .CI(n22975), .CO(n33089), .S(
        n22977) );
  AOI22XL U27744 ( .A0(n16657), .A1(n22977), .B0(conv_1[385]), .B1(n22976), 
        .Y(n22978) );
  NAND2XL U27745 ( .A(n22978), .B(n34696), .Y(n16078) );
  NAND2XL U27746 ( .A(n27632), .B(n34525), .Y(n28821) );
  AND2XL U27747 ( .A(n22982), .B(n22981), .Y(n23140) );
  INVXL U27748 ( .A(conv_1[335]), .Y(n22992) );
  AOI2BB1XL U27749 ( .A0N(conv_1[335]), .A1N(n22994), .B0(n28821), .Y(n22983)
         );
  AOI2BB1XL U27750 ( .A0N(n35434), .A1N(n22993), .B0(n22983), .Y(n22985) );
  NAND2XL U27751 ( .A(conv_1[336]), .B(n22985), .Y(n22984) );
  OAI211XL U27752 ( .A0(conv_1[336]), .A1(n22985), .B0(n27932), .C0(n22984), 
        .Y(n22986) );
  OAI211XL U27753 ( .A0(n35437), .A1(n22987), .B0(n34281), .C0(n22986), .Y(
        n16127) );
  AOI21XL U27754 ( .A0(n22994), .A1(n35434), .B0(n22988), .Y(n22990) );
  NAND2XL U27755 ( .A(conv_1[335]), .B(n22990), .Y(n22989) );
  OAI211XL U27756 ( .A0(conv_1[335]), .A1(n22990), .B0(n27932), .C0(n22989), 
        .Y(n22991) );
  OAI211XL U27757 ( .A0(n35437), .A1(n22992), .B0(n34682), .C0(n22991), .Y(
        n16128) );
  NAND2XL U27758 ( .A(conv_1[336]), .B(n22993), .Y(n22999) );
  OAI31XL U27759 ( .A0(conv_1[335]), .A1(conv_1[336]), .A2(n22994), .B0(n35434), .Y(n22998) );
  OAI2BB1XL U27760 ( .A0N(n28821), .A1N(n22999), .B0(n22998), .Y(n22996) );
  NAND2XL U27761 ( .A(n23000), .B(n22996), .Y(n22995) );
  OAI211XL U27762 ( .A0(n23000), .A1(n22996), .B0(n27932), .C0(n22995), .Y(
        n22997) );
  OAI211XL U27763 ( .A0(n35437), .A1(n23000), .B0(n34544), .C0(n22997), .Y(
        n16126) );
  INVXL U27764 ( .A(conv_1[341]), .Y(n28823) );
  AOI21XL U27765 ( .A0(n23000), .A1(n22998), .B0(n28821), .Y(n35432) );
  AOI2BB1XL U27766 ( .A0N(conv_1[339]), .A1N(n23010), .B0(n28821), .Y(n23004)
         );
  OAI21XL U27767 ( .A0(conv_1[340]), .A1(n23004), .B0(n35434), .Y(n28822) );
  NAND2XL U27768 ( .A(conv_1[338]), .B(n35433), .Y(n23011) );
  OAI2BB1XL U27769 ( .A0N(conv_1[340]), .A1N(n23005), .B0(n28821), .Y(n33884)
         );
  NAND2XL U27770 ( .A(n28822), .B(n33884), .Y(n23002) );
  NAND2XL U27771 ( .A(n28823), .B(n23002), .Y(n23001) );
  OAI211XL U27772 ( .A0(n28823), .A1(n23002), .B0(n33788), .C0(n23001), .Y(
        n23003) );
  OAI211XL U27773 ( .A0(n35437), .A1(n28823), .B0(n16652), .C0(n23003), .Y(
        n16122) );
  AOI2BB1XL U27774 ( .A0N(n35434), .A1N(n23005), .B0(n23004), .Y(n23007) );
  NAND2XL U27775 ( .A(conv_1[340]), .B(n23007), .Y(n23006) );
  OAI211XL U27776 ( .A0(conv_1[340]), .A1(n23007), .B0(n27932), .C0(n23006), 
        .Y(n23008) );
  OAI211XL U27777 ( .A0(n35437), .A1(n23009), .B0(n16652), .C0(n23008), .Y(
        n16123) );
  AOI21XL U27778 ( .A0(n28821), .A1(n23011), .B0(n23010), .Y(n23013) );
  NAND2XL U27779 ( .A(conv_1[339]), .B(n23013), .Y(n23012) );
  OAI211XL U27780 ( .A0(conv_1[339]), .A1(n23013), .B0(n27932), .C0(n23012), 
        .Y(n23014) );
  OAI211XL U27781 ( .A0(n35437), .A1(n23015), .B0(n34682), .C0(n23014), .Y(
        n16124) );
  AOI222XL U27782 ( .A0(n23016), .A1(n23278), .B0(n23781), .B1(n23276), .C0(
        n23784), .C1(n23272), .Y(n23285) );
  NAND2XL U27783 ( .A(conv_1[390]), .B(n30649), .Y(n30648) );
  OAI21XL U27784 ( .A0(n35272), .A1(n32016), .B0(n30648), .Y(n30667) );
  AOI21XL U27785 ( .A0(conv_1[391]), .A1(n30667), .B0(n30666), .Y(n30486) );
  NAND2XL U27786 ( .A(n24909), .B(n27990), .Y(n30485) );
  AND2XL U27787 ( .A(n30485), .B(n30486), .Y(n30487) );
  INVXL U27788 ( .A(conv_1[392]), .Y(n30492) );
  OAI22XL U27789 ( .A0(n30486), .A1(n30485), .B0(n30487), .B1(n30492), .Y(
        n27633) );
  AOI22XL U27790 ( .A0(n32181), .A1(n23021), .B0(conv_1[393]), .B1(n33649), 
        .Y(n23022) );
  NAND2XL U27791 ( .A(n23022), .B(n32867), .Y(n16070) );
  INVXL U27792 ( .A(conv_1[434]), .Y(n29334) );
  AOI22XL U27793 ( .A0(n33712), .A1(intadd_1_SUM_0_), .B0(conv_1[423]), .B1(
        n35510), .Y(n23023) );
  NAND2XL U27794 ( .A(n23023), .B(n32867), .Y(n16040) );
  NAND2XL U27795 ( .A(conv_2[45]), .B(n28124), .Y(n23024) );
  NAND2XL U27796 ( .A(n34506), .B(n28126), .Y(n23825) );
  AOI21XL U27797 ( .A0(n18913), .A1(n23024), .B0(n27799), .Y(n23826) );
  NAND2XL U27798 ( .A(conv_2[46]), .B(n23826), .Y(n23025) );
  NAND2XL U27799 ( .A(n23825), .B(n23025), .Y(n23027) );
  NAND2XL U27800 ( .A(n35853), .B(n23027), .Y(n23026) );
  NAND2XL U27801 ( .A(n23027), .B(n28128), .Y(n23028) );
  OAI2BB1XL U27802 ( .A0N(conv_2[47]), .A1N(n31067), .B0(n23028), .Y(n27800)
         );
  AOI22XL U27803 ( .A0(n32660), .A1(n23029), .B0(conv_2[48]), .B1(n30873), .Y(
        n23030) );
  NAND2XL U27804 ( .A(n23030), .B(n34105), .Y(n15272) );
  AOI22XL U27805 ( .A0(n32660), .A1(n23034), .B0(conv_2[93]), .B1(n23033), .Y(
        n23035) );
  NAND2XL U27806 ( .A(n23035), .B(n34105), .Y(n15269) );
  AOI22XL U27807 ( .A0(n32660), .A1(intadd_0_SUM_1_), .B0(conv_2[3]), .B1(
        n33566), .Y(n23036) );
  NAND2XL U27808 ( .A(n23036), .B(n34105), .Y(n15275) );
  AOI22XL U27809 ( .A0(n33712), .A1(n23039), .B0(conv_2[138]), .B1(n35909), 
        .Y(n23040) );
  NAND2XL U27810 ( .A(n23040), .B(n34105), .Y(n15266) );
  NAND2XL U27811 ( .A(conv_2[120]), .B(n28124), .Y(n23041) );
  NAND2XL U27812 ( .A(n34492), .B(n28126), .Y(n23847) );
  AOI21XL U27813 ( .A0(n18913), .A1(n23041), .B0(n28948), .Y(n23848) );
  NAND2XL U27814 ( .A(conv_2[121]), .B(n23848), .Y(n23042) );
  NAND2XL U27815 ( .A(n23847), .B(n23042), .Y(n23044) );
  NAND2XL U27816 ( .A(n35853), .B(n23044), .Y(n23043) );
  OAI31XL U27817 ( .A0(n35853), .A1(n28948), .A2(n23044), .B0(n23043), .Y(
        n30003) );
  NAND2XL U27818 ( .A(n23044), .B(n28128), .Y(n23045) );
  OAI2BB1XL U27819 ( .A0N(conv_2[122]), .A1N(n30003), .B0(n23045), .Y(n23333)
         );
  INVXL U27820 ( .A(conv_2[134]), .Y(n30448) );
  AOI22XL U27821 ( .A0(n32660), .A1(n23046), .B0(conv_2[123]), .B1(n33801), 
        .Y(n23047) );
  NAND2XL U27822 ( .A(n23047), .B(n34105), .Y(n15267) );
  AOI22XL U27823 ( .A0(n32660), .A1(n23050), .B0(conv_3[453]), .B1(n33774), 
        .Y(n23051) );
  NAND2XL U27824 ( .A(n23051), .B(n35574), .Y(n15785) );
  AOI22XL U27825 ( .A0(n25766), .A1(n23784), .B0(n34921), .B1(n23275), .Y(
        n23057) );
  OAI22XL U27826 ( .A0(n23282), .A1(n23053), .B0(n23789), .B1(n23052), .Y(
        n23054) );
  INVXL U27827 ( .A(conv_3[481]), .Y(n30529) );
  NAND2XL U27828 ( .A(conv_3[480]), .B(n29678), .Y(n23059) );
  OAI2BB1XL U27829 ( .A0N(n30536), .A1N(n23059), .B0(n33530), .Y(n30524) );
  NAND3XL U27830 ( .A(conv_3[480]), .B(n33530), .C(n29678), .Y(n31108) );
  OAI21XL U27831 ( .A0(n30529), .A1(n30524), .B0(n23060), .Y(n23061) );
  AOI21XL U27832 ( .A0(n33530), .A1(n27619), .B0(n23061), .Y(n30497) );
  INVXL U27833 ( .A(conv_3[482]), .Y(n30502) );
  NAND2XL U27834 ( .A(n27619), .B(n23061), .Y(n30498) );
  OAI21XL U27835 ( .A0(n30497), .A1(n30502), .B0(n30498), .Y(n23514) );
  INVXL U27836 ( .A(conv_3[494]), .Y(n32233) );
  AOI22XL U27837 ( .A0(n32660), .A1(n23062), .B0(conv_3[483]), .B1(n35833), 
        .Y(n23063) );
  NAND2XL U27838 ( .A(n23063), .B(n35574), .Y(n15783) );
  NAND2XL U27839 ( .A(conv_3[285]), .B(n30619), .Y(n30618) );
  OAI21XL U27840 ( .A0(n30536), .A1(n31871), .B0(n30618), .Y(n23064) );
  INVXL U27841 ( .A(n23064), .Y(n30537) );
  INVXL U27842 ( .A(conv_3[286]), .Y(n30542) );
  OAI22XL U27843 ( .A0(n30536), .A1(n30618), .B0(n30537), .B1(n30542), .Y(
        n31085) );
  INVXL U27844 ( .A(conv_3[299]), .Y(n32240) );
  AOI22XL U27845 ( .A0(n33712), .A1(n23067), .B0(conv_3[289]), .B1(n32566), 
        .Y(n23068) );
  NAND2XL U27846 ( .A(n23068), .B(n34097), .Y(n15760) );
  ADDFX1 U27847 ( .A(conv_3[379]), .B(n23070), .CI(n23069), .CO(n31455), .S(
        n23071) );
  AOI22XL U27848 ( .A0(n32660), .A1(n23071), .B0(conv_3[379]), .B1(n32623), 
        .Y(n23072) );
  NAND2XL U27849 ( .A(n23072), .B(n34097), .Y(n15754) );
  NAND2XL U27850 ( .A(n28068), .B(n27535), .Y(n23076) );
  NAND2XL U27851 ( .A(n23988), .B(conv_2[375]), .Y(n23987) );
  INVXL U27852 ( .A(n23987), .Y(n23073) );
  NAND2XL U27853 ( .A(n23073), .B(n28126), .Y(n23074) );
  OAI32XL U27854 ( .A0(n23073), .A1(n27532), .A2(n18913), .B0(n28126), .B1(
        n23987), .Y(n30299) );
  NAND2XL U27855 ( .A(n23074), .B(n30298), .Y(n30400) );
  NOR2X1 U27856 ( .A(conv_2[383]), .B(n33673), .Y(n33674) );
  NOR2X1 U27857 ( .A(n33674), .B(n36025), .Y(n28012) );
  NAND2XL U27858 ( .A(n33417), .B(conv_2[381]), .Y(n36024) );
  INVXL U27859 ( .A(conv_2[382]), .Y(n36027) );
  AOI22XL U27860 ( .A0(n16656), .A1(n23080), .B0(conv_2[385]), .B1(n34531), 
        .Y(n23081) );
  NAND2XL U27861 ( .A(n23081), .B(n35859), .Y(n14948) );
  NAND2XL U27862 ( .A(conv_2[330]), .B(n28124), .Y(n23082) );
  AOI21XL U27863 ( .A0(n18913), .A1(n23082), .B0(n34522), .Y(n29810) );
  NAND2XL U27864 ( .A(n34485), .B(n28126), .Y(n29809) );
  OAI2BB1XL U27865 ( .A0N(conv_2[331]), .A1N(n29810), .B0(n29809), .Y(n23084)
         );
  NAND2XL U27866 ( .A(n35853), .B(n23084), .Y(n23083) );
  OAI31XL U27867 ( .A0(n35853), .A1(n34522), .A2(n23084), .B0(n23083), .Y(
        n29999) );
  NAND2XL U27868 ( .A(n23084), .B(n28128), .Y(n23085) );
  OAI2BB1XL U27869 ( .A0N(conv_2[332]), .A1N(n29999), .B0(n23085), .Y(n24301)
         );
  AOI222XL U27870 ( .A0(conv_2[334]), .A1(n23867), .B0(conv_2[334]), .B1(
        n23868), .C0(n23867), .C1(n23868), .Y(n23086) );
  NAND2XL U27871 ( .A(n35997), .B(n23086), .Y(n28097) );
  OAI21XL U27872 ( .A0(conv_2[335]), .A1(n28096), .B0(n35995), .Y(n35989) );
  AOI22XL U27873 ( .A0(n16657), .A1(n23087), .B0(conv_2[337]), .B1(n24303), 
        .Y(n23088) );
  NAND2XL U27874 ( .A(n23088), .B(n35859), .Y(n14981) );
  INVXL U27875 ( .A(conv_2[345]), .Y(n34418) );
  NAND2XL U27876 ( .A(n23096), .B(n34762), .Y(n34416) );
  INVXL U27877 ( .A(conv_2[346]), .Y(n24490) );
  INVXL U27878 ( .A(n23097), .Y(n23095) );
  OAI211XL U27879 ( .A0(n23096), .A1(n28126), .B0(n34762), .C0(n23095), .Y(
        n24488) );
  OAI21XL U27880 ( .A0(n35853), .A1(n26717), .B0(n29878), .Y(n23098) );
  INVXL U27881 ( .A(n23098), .Y(n29879) );
  INVXL U27882 ( .A(conv_2[347]), .Y(n29884) );
  OAI22XL U27883 ( .A0(n35853), .A1(n29878), .B0(n29879), .B1(n29884), .Y(
        n23712) );
  INVXL U27884 ( .A(conv_2[350]), .Y(n33931) );
  AOI22XL U27885 ( .A0(n34028), .A1(n23099), .B0(conv_2[351]), .B1(n24190), 
        .Y(n23100) );
  NAND2XL U27886 ( .A(n23100), .B(n35859), .Y(n14972) );
  INVXL U27887 ( .A(n22269), .Y(n34465) );
  NAND3XL U27888 ( .A(n34465), .B(conv_2[315]), .C(n28124), .Y(n23101) );
  INVXL U27889 ( .A(conv_2[316]), .Y(n23459) );
  INVXL U27890 ( .A(n23101), .Y(n34463) );
  AOI32XL U27891 ( .A0(n34465), .A1(n28126), .A2(n23101), .B0(n34463), .B1(
        n18913), .Y(n23457) );
  NOR2X1 U27892 ( .A(n23459), .B(n23457), .Y(n23455) );
  AOI21XL U27893 ( .A0(n34465), .A1(n28128), .B0(n23103), .Y(n29872) );
  INVXL U27894 ( .A(conv_2[317]), .Y(n29877) );
  NAND2XL U27895 ( .A(n28128), .B(n23103), .Y(n29873) );
  NOR2X1 U27896 ( .A(n23105), .B(n23104), .Y(n28865) );
  NOR2X1 U27897 ( .A(n35982), .B(n23106), .Y(n28051) );
  AOI22XL U27898 ( .A0(n32181), .A1(n23107), .B0(conv_2[321]), .B1(n24298), 
        .Y(n23108) );
  NAND2XL U27899 ( .A(n23108), .B(n35859), .Y(n14992) );
  NAND2XL U27900 ( .A(n29046), .B(n34579), .Y(n23115) );
  NAND2XL U27901 ( .A(conv_2[150]), .B(n28124), .Y(n23109) );
  AOI221XL U27902 ( .A0(n34578), .A1(n28126), .B0(n23109), .B1(n18913), .C0(
        n23296), .Y(n23863) );
  NAND2XL U27903 ( .A(n34578), .B(n28126), .Y(n23110) );
  OAI2BB1XL U27904 ( .A0N(conv_2[151]), .A1N(n23863), .B0(n23110), .Y(n24255)
         );
  AND2XL U27905 ( .A(n23112), .B(n23111), .Y(n23266) );
  INVXL U27906 ( .A(n23267), .Y(n23113) );
  OAI21XL U27907 ( .A0(conv_2[153]), .A1(n23266), .B0(n23113), .Y(n23114) );
  AOI22XL U27908 ( .A0(n33157), .A1(n23116), .B0(conv_2[156]), .B1(n24358), 
        .Y(n23117) );
  NAND2XL U27909 ( .A(n23117), .B(n35859), .Y(n15102) );
  NAND2XL U27910 ( .A(n29046), .B(n34502), .Y(n23124) );
  NAND3XL U27911 ( .A(n28124), .B(n34502), .C(conv_2[360]), .Y(n23118) );
  INVXL U27912 ( .A(n23118), .Y(n34501) );
  NAND2XL U27913 ( .A(n34501), .B(n28126), .Y(n23119) );
  OAI32XL U27914 ( .A0(n34501), .A1(n23504), .A2(n18913), .B0(n28126), .B1(
        n23118), .Y(n29806) );
  NAND2XL U27915 ( .A(n29806), .B(conv_2[361]), .Y(n29805) );
  NAND2XL U27916 ( .A(n23119), .B(n29805), .Y(n23121) );
  NAND2XL U27917 ( .A(n28128), .B(n23121), .Y(n23122) );
  NAND2XL U27918 ( .A(n35853), .B(n23121), .Y(n23120) );
  OAI31XL U27919 ( .A0(n35853), .A1(n23504), .A2(n23121), .B0(n23120), .Y(
        n29989) );
  NAND2XL U27920 ( .A(n29989), .B(conv_2[362]), .Y(n29988) );
  AOI222XL U27921 ( .A0(n23234), .A1(conv_2[363]), .B0(n23234), .B1(n23233), 
        .C0(conv_2[363]), .C1(n23233), .Y(n23123) );
  NAND2XL U27922 ( .A(n23124), .B(n23123), .Y(n23357) );
  NAND2XL U27923 ( .A(n27273), .B(n23125), .Y(n34564) );
  AOI21XL U27924 ( .A0(conv_2[368]), .A1(n29507), .B0(n34570), .Y(n29493) );
  INVXL U27925 ( .A(conv_2[374]), .Y(n29472) );
  AOI22XL U27926 ( .A0(n16657), .A1(n23126), .B0(conv_2[370]), .B1(n24455), 
        .Y(n23127) );
  NAND2XL U27927 ( .A(n23127), .B(n35859), .Y(n14958) );
  AOI21XL U27928 ( .A0(n33088), .A1(n23129), .B0(n23128), .Y(n23131) );
  NAND2XL U27929 ( .A(conv_1[382]), .B(n23131), .Y(n23130) );
  OAI211XL U27930 ( .A0(conv_1[382]), .A1(n23131), .B0(n24378), .C0(n23130), 
        .Y(n23132) );
  OAI211XL U27931 ( .A0(n35466), .A1(n23133), .B0(n16652), .C0(n23132), .Y(
        n16081) );
  AOI2BB1XL U27932 ( .A0N(n35463), .A1N(n23135), .B0(n23134), .Y(n23137) );
  NAND2XL U27933 ( .A(conv_1[381]), .B(n23137), .Y(n23136) );
  OAI211XL U27934 ( .A0(conv_1[381]), .A1(n23137), .B0(n33788), .C0(n23136), 
        .Y(n23138) );
  OAI211XL U27935 ( .A0(n35466), .A1(n23139), .B0(n34544), .C0(n23138), .Y(
        n16082) );
  INVXL U27936 ( .A(conv_1[333]), .Y(n23145) );
  NAND2XL U27937 ( .A(conv_1[333]), .B(n23143), .Y(n23142) );
  OAI211XL U27938 ( .A0(conv_1[333]), .A1(n23143), .B0(n27932), .C0(n23142), 
        .Y(n23144) );
  OAI211XL U27939 ( .A0(n35437), .A1(n23145), .B0(n23144), .C0(n32867), .Y(
        n16130) );
  INVXL U27940 ( .A(conv_2[240]), .Y(n23148) );
  NAND2XL U27941 ( .A(conv_2[240]), .B(n23146), .Y(n29768) );
  OAI211XL U27942 ( .A0(conv_2[240]), .A1(n23146), .B0(n30090), .C0(n29768), 
        .Y(n23147) );
  OAI211XL U27943 ( .A0(n35945), .A1(n23148), .B0(n23147), .C0(n34583), .Y(
        n15367) );
  NAND2XL U27944 ( .A(conv_1[370]), .B(n23153), .Y(n23152) );
  OAI211XL U27945 ( .A0(conv_1[370]), .A1(n23153), .B0(n32052), .C0(n23152), 
        .Y(n23154) );
  OAI211XL U27946 ( .A0(n35458), .A1(n23155), .B0(n16652), .C0(n23154), .Y(
        n16093) );
  OAI21XL U27947 ( .A0(n18913), .A1(n24021), .B0(n29768), .Y(n23156) );
  INVXL U27948 ( .A(n23156), .Y(n29769) );
  INVXL U27949 ( .A(conv_2[241]), .Y(n29774) );
  OAI22XL U27950 ( .A0(n18913), .A1(n29768), .B0(n29769), .B1(n29774), .Y(
        n30272) );
  AOI21XL U27951 ( .A0(n28145), .A1(n28146), .B0(n23157), .Y(n23159) );
  NAND2XL U27952 ( .A(conv_2[243]), .B(n23159), .Y(n23158) );
  OAI211XL U27953 ( .A0(conv_2[243]), .A1(n23159), .B0(n35336), .C0(n23158), 
        .Y(n23160) );
  OAI211XL U27954 ( .A0(n35945), .A1(n23161), .B0(n34105), .C0(n23160), .Y(
        n15259) );
  NAND2XL U27955 ( .A(n23164), .B(n23163), .Y(n23166) );
  NAND2XL U27956 ( .A(conv_1[298]), .B(n23166), .Y(n23165) );
  OAI211XL U27957 ( .A0(conv_1[298]), .A1(n23166), .B0(n24378), .C0(n23165), 
        .Y(n23167) );
  OAI211XL U27958 ( .A0(n34325), .A1(n23168), .B0(n16652), .C0(n23167), .Y(
        n16165) );
  INVXL U27959 ( .A(conv_1[292]), .Y(n23174) );
  NAND2XL U27960 ( .A(conv_1[292]), .B(n23172), .Y(n23171) );
  OAI211XL U27961 ( .A0(conv_1[292]), .A1(n23172), .B0(n27932), .C0(n23171), 
        .Y(n23173) );
  OAI211XL U27962 ( .A0(n34325), .A1(n23174), .B0(n16652), .C0(n23173), .Y(
        n16171) );
  OAI21XL U27963 ( .A0(n34319), .A1(n23176), .B0(n23175), .Y(n23178) );
  NAND2XL U27964 ( .A(n23180), .B(n23178), .Y(n23177) );
  OAI211XL U27965 ( .A0(n23180), .A1(n23178), .B0(n16657), .C0(n23177), .Y(
        n23179) );
  OAI211XL U27966 ( .A0(n34325), .A1(n23180), .B0(n34689), .C0(n23179), .Y(
        n16170) );
  AOI21XL U27967 ( .A0(n34319), .A1(n23182), .B0(n23181), .Y(n23184) );
  NAND2XL U27968 ( .A(conv_1[294]), .B(n23184), .Y(n23183) );
  OAI211XL U27969 ( .A0(conv_1[294]), .A1(n23184), .B0(n30090), .C0(n23183), 
        .Y(n23185) );
  OAI211XL U27970 ( .A0(n34325), .A1(n23186), .B0(n34689), .C0(n23185), .Y(
        n16169) );
  INVXL U27971 ( .A(conv_1[295]), .Y(n23192) );
  AOI2BB1XL U27972 ( .A0N(n34319), .A1N(n23188), .B0(n23187), .Y(n23190) );
  NAND2XL U27973 ( .A(conv_1[295]), .B(n23190), .Y(n23189) );
  OAI211XL U27974 ( .A0(conv_1[295]), .A1(n23190), .B0(n32052), .C0(n23189), 
        .Y(n23191) );
  OAI211XL U27975 ( .A0(n34325), .A1(n23192), .B0(n34689), .C0(n23191), .Y(
        n16168) );
  INVXL U27976 ( .A(conv_1[378]), .Y(n23198) );
  XOR2XL U27977 ( .A(n23194), .B(n23193), .Y(n23196) );
  NAND2XL U27978 ( .A(conv_1[378]), .B(n23196), .Y(n23195) );
  OAI211XL U27979 ( .A0(conv_1[378]), .A1(n23196), .B0(n33778), .C0(n23195), 
        .Y(n23197) );
  OAI211XL U27980 ( .A0(n35466), .A1(n23198), .B0(n32867), .C0(n23197), .Y(
        n16085) );
  NAND2XL U27981 ( .A(n29680), .B(n34507), .Y(n23199) );
  NAND2XL U27982 ( .A(n30536), .B(n23201), .Y(n23200) );
  OAI211XL U27983 ( .A0(n30536), .A1(n23201), .B0(n34507), .C0(n23200), .Y(
        n23744) );
  INVXL U27984 ( .A(conv_3[46]), .Y(n23746) );
  OAI21XL U27985 ( .A0(n18997), .A1(n27799), .B0(n23203), .Y(n23204) );
  INVXL U27986 ( .A(n23204), .Y(n30748) );
  AOI222XL U27987 ( .A0(n29720), .A1(n29719), .B0(n29720), .B1(conv_3[48]), 
        .C0(n29719), .C1(conv_3[48]), .Y(n23205) );
  INVXL U27988 ( .A(n23205), .Y(n23207) );
  NAND2XL U27989 ( .A(n23207), .B(n23206), .Y(n23928) );
  OR2XL U27990 ( .A(n23207), .B(n23206), .Y(n23929) );
  AND2XL U27991 ( .A(n23928), .B(n23929), .Y(n23209) );
  NAND2XL U27992 ( .A(conv_3[49]), .B(n23209), .Y(n23208) );
  OAI211XL U27993 ( .A0(conv_3[49]), .A1(n23209), .B0(n35336), .C0(n23208), 
        .Y(n23210) );
  OAI211XL U27994 ( .A0(n34392), .A1(n23211), .B0(n34097), .C0(n23210), .Y(
        n15776) );
  INVXL U27995 ( .A(conv_2[404]), .Y(n33262) );
  INVXL U27996 ( .A(conv_2[390]), .Y(n23214) );
  NAND2XL U27997 ( .A(n23212), .B(conv_2[390]), .Y(n24445) );
  OAI211XL U27998 ( .A0(n23212), .A1(conv_2[390]), .B0(n30090), .C0(n24445), 
        .Y(n23213) );
  OAI211XL U27999 ( .A0(n36031), .A1(n23214), .B0(n34583), .C0(n23213), .Y(
        n15357) );
  INVXL U28000 ( .A(conv_3[314]), .Y(n33115) );
  NAND2XL U28001 ( .A(conv_3[300]), .B(n29678), .Y(n23216) );
  NAND2XL U28002 ( .A(n27058), .B(n29680), .Y(n23217) );
  INVXL U28003 ( .A(n23217), .Y(n23215) );
  NAND2XL U28004 ( .A(n31023), .B(conv_3[301]), .Y(n31022) );
  NAND2XL U28005 ( .A(n23217), .B(n31022), .Y(n23218) );
  NAND2XL U28006 ( .A(n27619), .B(n23218), .Y(n30714) );
  NAND2XL U28007 ( .A(conv_3[302]), .B(n30713), .Y(n23220) );
  AOI222XL U28008 ( .A0(n23486), .A1(conv_3[303]), .B0(n23486), .B1(n23485), 
        .C0(conv_3[303]), .C1(n23485), .Y(n23221) );
  INVXL U28009 ( .A(n23221), .Y(n23222) );
  NOR2X1 U28010 ( .A(n23223), .B(n23222), .Y(n31404) );
  NAND2XL U28011 ( .A(conv_3[304]), .B(n23225), .Y(n23224) );
  OAI211XL U28012 ( .A0(conv_3[304]), .A1(n23225), .B0(n33822), .C0(n23224), 
        .Y(n23226) );
  OAI211XL U28013 ( .A0(n35736), .A1(n23227), .B0(n34097), .C0(n23226), .Y(
        n15759) );
  INVXL U28014 ( .A(conv_2[106]), .Y(n23572) );
  OAI21XL U28015 ( .A0(n18913), .A1(n34715), .B0(n23574), .Y(n23228) );
  INVXL U28016 ( .A(n23228), .Y(n23573) );
  NAND2XL U28017 ( .A(conv_2[106]), .B(n23231), .Y(n23230) );
  OAI211XL U28018 ( .A0(conv_2[106]), .A1(n23231), .B0(n33982), .C0(n23230), 
        .Y(n23232) );
  OAI211XL U28019 ( .A0(n35894), .A1(n23572), .B0(n23232), .C0(n35847), .Y(
        n15340) );
  INVXL U28020 ( .A(conv_2[363]), .Y(n23238) );
  NAND2XL U28021 ( .A(conv_2[363]), .B(n23236), .Y(n23235) );
  OAI211XL U28022 ( .A0(conv_2[363]), .A1(n23236), .B0(n33822), .C0(n23235), 
        .Y(n23237) );
  OAI211XL U28023 ( .A0(n36017), .A1(n23238), .B0(n23237), .C0(n34105), .Y(
        n15251) );
  INVXL U28024 ( .A(conv_2[510]), .Y(n23255) );
  AOI22XL U28025 ( .A0(n18197), .A1(n23240), .B0(n18463), .B1(n23239), .Y(
        n23251) );
  AOI22XL U28026 ( .A0(n28324), .A1(n23242), .B0(n26376), .B1(n23241), .Y(
        n23246) );
  AOI22XL U28027 ( .A0(n26262), .A1(n23244), .B0(n16670), .B1(n23243), .Y(
        n23245) );
  OAI211XL U28028 ( .A0(conv_2[510]), .A1(n23253), .B0(n33982), .C0(n23565), 
        .Y(n23254) );
  OAI211XL U28029 ( .A0(n31013), .A1(n23255), .B0(n23254), .C0(n34583), .Y(
        n15349) );
  INVXL U28030 ( .A(conv_3[524]), .Y(n31296) );
  INVXL U28031 ( .A(conv_3[514]), .Y(n23265) );
  NAND2XL U28032 ( .A(conv_3[510]), .B(n29678), .Y(n23256) );
  AOI21XL U28033 ( .A0(n30536), .A1(n23256), .B0(n27764), .Y(n30519) );
  NAND2XL U28034 ( .A(n27062), .B(n29680), .Y(n30518) );
  OAI2BB1XL U28035 ( .A0N(conv_3[511]), .A1N(n30519), .B0(n30518), .Y(n23258)
         );
  NAND2XL U28036 ( .A(n18997), .B(n23258), .Y(n23257) );
  OAI31XL U28037 ( .A0(n18997), .A1(n27764), .A2(n23258), .B0(n23257), .Y(
        n30720) );
  NAND2XL U28038 ( .A(n23258), .B(n27619), .Y(n23259) );
  OAI2BB1XL U28039 ( .A0N(conv_3[512]), .A1N(n30720), .B0(n23259), .Y(n23738)
         );
  AND2XL U28040 ( .A(n23261), .B(n23260), .Y(n24459) );
  NAND2XL U28041 ( .A(conv_3[514]), .B(n23263), .Y(n23262) );
  OAI211XL U28042 ( .A0(conv_3[514]), .A1(n23263), .B0(n35336), .C0(n23262), 
        .Y(n23264) );
  OAI211XL U28043 ( .A0(n33303), .A1(n23265), .B0(n34097), .C0(n23264), .Y(
        n15745) );
  INVXL U28044 ( .A(conv_2[153]), .Y(n23271) );
  NAND2XL U28045 ( .A(conv_2[153]), .B(n23269), .Y(n23268) );
  OAI211XL U28046 ( .A0(conv_2[153]), .A1(n23269), .B0(n35336), .C0(n23268), 
        .Y(n23270) );
  OAI211XL U28047 ( .A0(n34631), .A1(n23271), .B0(n23270), .C0(n34105), .Y(
        n15265) );
  NAND2XL U28048 ( .A(n23274), .B(n23782), .Y(n23284) );
  INVXL U28049 ( .A(n23272), .Y(n23281) );
  AOI22XL U28050 ( .A0(n23276), .A1(n23275), .B0(n23274), .B1(n23273), .Y(
        n23280) );
  NAND2XL U28051 ( .A(n23278), .B(n23277), .Y(n23279) );
  INVXL U28052 ( .A(n23786), .Y(n23283) );
  NAND2XL U28053 ( .A(conv_1[210]), .B(n30672), .Y(n23286) );
  NAND2XL U28054 ( .A(n33869), .B(n27429), .Y(n33030) );
  AOI21XL U28055 ( .A0(n35272), .A1(n23286), .B0(n28660), .Y(n33031) );
  NAND2XL U28056 ( .A(conv_1[211]), .B(n33031), .Y(n33028) );
  NAND2XL U28057 ( .A(n33030), .B(n33028), .Y(n23288) );
  NAND2XL U28058 ( .A(n33403), .B(n23288), .Y(n23287) );
  OAI31XL U28059 ( .A0(n33403), .A1(n28660), .A2(n23288), .B0(n23287), .Y(
        n23906) );
  NAND2XL U28060 ( .A(n23288), .B(n24909), .Y(n23289) );
  OAI2BB1XL U28061 ( .A0N(conv_1[212]), .A1N(n23906), .B0(n23289), .Y(n24291)
         );
  AOI222XL U28062 ( .A0(n23998), .A1(n23999), .B0(n23998), .B1(conv_1[214]), 
        .C0(n23999), .C1(conv_1[214]), .Y(n23290) );
  OAI21XL U28063 ( .A0(conv_1[217]), .A1(n35390), .B0(n35392), .Y(n24680) );
  NAND2XL U28064 ( .A(n24684), .B(n24680), .Y(n23291) );
  NAND2XL U28065 ( .A(n35392), .B(n23291), .Y(n34538) );
  NAND2XL U28066 ( .A(n34543), .B(n34538), .Y(n25437) );
  NAND2XL U28067 ( .A(n28602), .B(n23290), .Y(n23342) );
  NAND2XL U28068 ( .A(conv_1[215]), .B(n23342), .Y(n23304) );
  OAI2BB1XL U28069 ( .A0N(conv_1[217]), .A1N(n35391), .B0(n28602), .Y(n24679)
         );
  AND2XL U28070 ( .A(n23291), .B(n24679), .Y(n34539) );
  OAI2BB1XL U28071 ( .A0N(conv_1[219]), .A1N(n34539), .B0(n28602), .Y(n25438)
         );
  OAI2BB1XL U28072 ( .A0N(n35392), .A1N(n25437), .B0(n25438), .Y(n23293) );
  NAND2XL U28073 ( .A(n23295), .B(n23293), .Y(n23292) );
  OAI211XL U28074 ( .A0(n23295), .A1(n23293), .B0(n33157), .C0(n23292), .Y(
        n23294) );
  OAI211XL U28075 ( .A0(n35395), .A1(n23295), .B0(n16652), .C0(n23294), .Y(
        n16243) );
  NAND2XL U28076 ( .A(conv_1[150]), .B(n26691), .Y(n26690) );
  INVXL U28077 ( .A(n26690), .Y(n23297) );
  AOI21XL U28078 ( .A0(n27429), .A1(n34579), .B0(n23297), .Y(n32794) );
  INVXL U28079 ( .A(conv_1[151]), .Y(n32799) );
  NAND2XL U28080 ( .A(n27429), .B(n23297), .Y(n32795) );
  OAI21XL U28081 ( .A0(n32794), .A1(n32799), .B0(n32795), .Y(n24427) );
  AOI222XL U28082 ( .A0(conv_1[154]), .A1(n24008), .B0(conv_1[154]), .B1(
        n24009), .C0(n24008), .C1(n24009), .Y(n23298) );
  INVXL U28083 ( .A(conv_1[155]), .Y(n23404) );
  NAND2XL U28084 ( .A(conv_1[158]), .B(n34043), .Y(n23393) );
  OAI2BB1XL U28085 ( .A0N(conv_1[160]), .A1N(n23388), .B0(n23394), .Y(n23381)
         );
  NAND4XL U28086 ( .A(conv_1[161]), .B(conv_1[162]), .C(n23394), .D(n23381), 
        .Y(n23412) );
  INVXL U28087 ( .A(conv_1[162]), .Y(n23380) );
  INVXL U28088 ( .A(conv_1[161]), .Y(n23386) );
  OAI31XL U28089 ( .A0(conv_1[158]), .A1(conv_1[159]), .A2(n34043), .B0(n34044), .Y(n23387) );
  OAI2BB1XL U28090 ( .A0N(n23392), .A1N(n23387), .B0(n34044), .Y(n23382) );
  NAND2XL U28091 ( .A(n23386), .B(n23382), .Y(n23299) );
  NAND3XL U28092 ( .A(n34044), .B(n23380), .C(n23376), .Y(n23411) );
  INVXL U28093 ( .A(conv_1[163]), .Y(n23416) );
  AOI22XL U28094 ( .A0(conv_1[163]), .A1(n23412), .B0(n23411), .B1(n23416), 
        .Y(n23301) );
  NAND2XL U28095 ( .A(conv_1[164]), .B(n23301), .Y(n23300) );
  OAI211XL U28096 ( .A0(conv_1[164]), .A1(n23301), .B0(n24499), .C0(n23300), 
        .Y(n23302) );
  OAI211XL U28097 ( .A0(n34676), .A1(n23375), .B0(n34696), .C0(n23302), .Y(
        n16299) );
  AOI21XL U28098 ( .A0(n28602), .A1(n23304), .B0(n23303), .Y(n23306) );
  NAND2XL U28099 ( .A(conv_1[216]), .B(n23306), .Y(n23305) );
  OAI211XL U28100 ( .A0(conv_1[216]), .A1(n23306), .B0(n24378), .C0(n23305), 
        .Y(n23307) );
  OAI211XL U28101 ( .A0(n35395), .A1(n23308), .B0(n16652), .C0(n23307), .Y(
        n16247) );
  NAND2XL U28102 ( .A(conv_1[324]), .B(n23312), .Y(n23311) );
  OAI211XL U28103 ( .A0(conv_1[324]), .A1(n23312), .B0(n27932), .C0(n23311), 
        .Y(n23313) );
  OAI211XL U28104 ( .A0(n34263), .A1(n23314), .B0(n34682), .C0(n23313), .Y(
        n16139) );
  AOI2BB1XL U28105 ( .A0N(n34259), .A1N(n23316), .B0(n23315), .Y(n23318) );
  NAND2XL U28106 ( .A(conv_1[323]), .B(n23318), .Y(n23317) );
  OAI211XL U28107 ( .A0(conv_1[323]), .A1(n23318), .B0(n27932), .C0(n23317), 
        .Y(n23319) );
  OAI211XL U28108 ( .A0(n34263), .A1(n23320), .B0(n16652), .C0(n23319), .Y(
        n16140) );
  OAI2BB1XL U28109 ( .A0N(n29382), .A1N(n23322), .B0(n23321), .Y(n23324) );
  NAND2XL U28110 ( .A(n23326), .B(n23324), .Y(n23323) );
  OAI211XL U28111 ( .A0(n23326), .A1(n23324), .B0(n27932), .C0(n23323), .Y(
        n23325) );
  OAI211XL U28112 ( .A0(n34263), .A1(n23326), .B0(n34689), .C0(n23325), .Y(
        n16141) );
  NAND2XL U28113 ( .A(n23328), .B(n23327), .Y(n23330) );
  NAND2XL U28114 ( .A(conv_1[328]), .B(n23330), .Y(n23329) );
  OAI211XL U28115 ( .A0(conv_1[328]), .A1(n23330), .B0(n27932), .C0(n23329), 
        .Y(n23331) );
  OAI211XL U28116 ( .A0(n34263), .A1(n23332), .B0(n34696), .C0(n23331), .Y(
        n16135) );
  INVXL U28117 ( .A(conv_2[124]), .Y(n23340) );
  NAND2XL U28118 ( .A(conv_2[124]), .B(n23338), .Y(n23337) );
  OAI211XL U28119 ( .A0(conv_2[124]), .A1(n23338), .B0(n32052), .C0(n23337), 
        .Y(n23339) );
  OAI211XL U28120 ( .A0(n34491), .A1(n23340), .B0(n34408), .C0(n23339), .Y(
        n15231) );
  INVXL U28121 ( .A(conv_1[215]), .Y(n23346) );
  NOR2BXL U28122 ( .AN(n23342), .B(n23341), .Y(n23344) );
  NAND2XL U28123 ( .A(conv_1[215]), .B(n23344), .Y(n23343) );
  OAI211XL U28124 ( .A0(conv_1[215]), .A1(n23344), .B0(n24499), .C0(n23343), 
        .Y(n23345) );
  OAI211XL U28125 ( .A0(n35395), .A1(n23346), .B0(n16652), .C0(n23345), .Y(
        n16248) );
  INVXL U28126 ( .A(conv_2[179]), .Y(n34598) );
  INVXL U28127 ( .A(conv_2[168]), .Y(n23355) );
  INVXL U28128 ( .A(conv_2[165]), .Y(n34434) );
  NAND2XL U28129 ( .A(n34431), .B(n28126), .Y(n23348) );
  INVXL U28130 ( .A(n34431), .Y(n23347) );
  NAND2XL U28131 ( .A(n31091), .B(conv_2[166]), .Y(n31090) );
  NAND2XL U28132 ( .A(n28128), .B(n23350), .Y(n23351) );
  XOR2XL U28133 ( .A(n29002), .B(n29001), .Y(n23353) );
  NAND2XL U28134 ( .A(conv_2[168]), .B(n23353), .Y(n23352) );
  OAI211XL U28135 ( .A0(conv_2[168]), .A1(n23353), .B0(n27932), .C0(n23352), 
        .Y(n23354) );
  OAI211XL U28136 ( .A0(n34589), .A1(n23355), .B0(n34105), .C0(n23354), .Y(
        n15264) );
  INVXL U28137 ( .A(conv_2[364]), .Y(n23361) );
  NOR2BXL U28138 ( .AN(n23357), .B(n23356), .Y(n23359) );
  NAND2XL U28139 ( .A(conv_2[364]), .B(n23359), .Y(n23358) );
  OAI211XL U28140 ( .A0(conv_2[364]), .A1(n23359), .B0(n32656), .C0(n23358), 
        .Y(n23360) );
  OAI211XL U28141 ( .A0(n36017), .A1(n23361), .B0(n23360), .C0(n34408), .Y(
        n15215) );
  XOR2XL U28142 ( .A(n23364), .B(n23363), .Y(n23366) );
  NAND2XL U28143 ( .A(conv_1[228]), .B(n23366), .Y(n23365) );
  OAI211XL U28144 ( .A0(conv_1[228]), .A1(n23366), .B0(n32656), .C0(n23365), 
        .Y(n23367) );
  OAI211XL U28145 ( .A0(n35408), .A1(n23368), .B0(n23367), .C0(n32867), .Y(
        n16235) );
  INVXL U28146 ( .A(conv_2[154]), .Y(n23374) );
  NAND2XL U28147 ( .A(conv_2[154]), .B(n23372), .Y(n23371) );
  OAI211XL U28148 ( .A0(conv_2[154]), .A1(n23372), .B0(n32052), .C0(n23371), 
        .Y(n23373) );
  OAI211XL U28149 ( .A0(n34631), .A1(n23374), .B0(n34408), .C0(n23373), .Y(
        n15229) );
  AOI32XL U28150 ( .A0(conv_1[161]), .A1(n23376), .A2(n23381), .B0(n34044), 
        .B1(n23376), .Y(n23378) );
  NAND2XL U28151 ( .A(n23380), .B(n23378), .Y(n23377) );
  OAI211XL U28152 ( .A0(n23380), .A1(n23378), .B0(n24499), .C0(n23377), .Y(
        n23379) );
  OAI211XL U28153 ( .A0(n34048), .A1(n23380), .B0(n34682), .C0(n23379), .Y(
        n16301) );
  NAND2XL U28154 ( .A(n23382), .B(n23381), .Y(n23384) );
  NAND2XL U28155 ( .A(n23386), .B(n23384), .Y(n23383) );
  OAI211XL U28156 ( .A0(n23386), .A1(n23384), .B0(n24499), .C0(n23383), .Y(
        n23385) );
  OAI211XL U28157 ( .A0(n34048), .A1(n23386), .B0(n34682), .C0(n23385), .Y(
        n16302) );
  OAI21XL U28158 ( .A0(n34044), .A1(n23388), .B0(n23387), .Y(n23390) );
  NAND2XL U28159 ( .A(n23392), .B(n23390), .Y(n23389) );
  OAI211XL U28160 ( .A0(n23392), .A1(n23390), .B0(n24499), .C0(n23389), .Y(
        n23391) );
  OAI211XL U28161 ( .A0(n34048), .A1(n23392), .B0(n34544), .C0(n23391), .Y(
        n16303) );
  OAI32XL U28162 ( .A0(n23394), .A1(conv_1[158]), .A2(n34043), .B0(n34044), 
        .B1(n23393), .Y(n23396) );
  NAND2XL U28163 ( .A(conv_1[159]), .B(n23396), .Y(n23395) );
  OAI211XL U28164 ( .A0(conv_1[159]), .A1(n23396), .B0(n24499), .C0(n23395), 
        .Y(n23397) );
  OAI211XL U28165 ( .A0(n34048), .A1(n23398), .B0(n34281), .C0(n23397), .Y(
        n16304) );
  NAND2XL U28166 ( .A(conv_1[155]), .B(n23402), .Y(n23401) );
  OAI211XL U28167 ( .A0(conv_1[155]), .A1(n23402), .B0(n24499), .C0(n23401), 
        .Y(n23403) );
  OAI211XL U28168 ( .A0(n34048), .A1(n23404), .B0(n34696), .C0(n23403), .Y(
        n16308) );
  INVXL U28169 ( .A(conv_1[156]), .Y(n23410) );
  NAND2XL U28170 ( .A(conv_1[156]), .B(n23408), .Y(n23407) );
  OAI211XL U28171 ( .A0(conv_1[156]), .A1(n23408), .B0(n24499), .C0(n23407), 
        .Y(n23409) );
  OAI211XL U28172 ( .A0(n34048), .A1(n23410), .B0(n16652), .C0(n23409), .Y(
        n16307) );
  NAND2XL U28173 ( .A(n23412), .B(n23411), .Y(n23414) );
  NAND2XL U28174 ( .A(conv_1[163]), .B(n23414), .Y(n23413) );
  OAI211XL U28175 ( .A0(conv_1[163]), .A1(n23414), .B0(n24499), .C0(n23413), 
        .Y(n23415) );
  OAI211XL U28176 ( .A0(n34048), .A1(n23416), .B0(n34281), .C0(n23415), .Y(
        n16300) );
  INVXL U28177 ( .A(conv_1[509]), .Y(n27190) );
  INVXL U28178 ( .A(conv_1[503]), .Y(n23432) );
  NAND2XL U28179 ( .A(n27230), .B(n33424), .Y(n23426) );
  NAND2XL U28180 ( .A(n27429), .B(n33424), .Y(n23417) );
  NAND2XL U28181 ( .A(conv_1[495]), .B(n30672), .Y(n33421) );
  NAND2XL U28182 ( .A(n35272), .B(n33421), .Y(n23418) );
  OAI211XL U28183 ( .A0(n35272), .A1(n33421), .B0(n33424), .C0(n23418), .Y(
        n24945) );
  INVXL U28184 ( .A(conv_1[496]), .Y(n24947) );
  OAI21XL U28185 ( .A0(n33403), .A1(n33422), .B0(n23420), .Y(n27474) );
  OR2XL U28186 ( .A(n33403), .B(n23420), .Y(n27472) );
  NAND2XL U28187 ( .A(n23421), .B(n27472), .Y(n27473) );
  AND2XL U28188 ( .A(n27474), .B(n27473), .Y(n23422) );
  AND2XL U28189 ( .A(n23423), .B(n23422), .Y(n29541) );
  INVXL U28190 ( .A(n29542), .Y(n23424) );
  OAI21XL U28191 ( .A0(conv_1[498]), .A1(n29541), .B0(n23424), .Y(n23425) );
  AND2XL U28192 ( .A(n23426), .B(n23425), .Y(n30696) );
  NAND2XL U28193 ( .A(n27131), .B(n26335), .Y(n26334) );
  AOI21XL U28194 ( .A0(n27119), .A1(n27131), .B0(n23428), .Y(n23430) );
  NAND2XL U28195 ( .A(conv_1[503]), .B(n23430), .Y(n23429) );
  OAI211XL U28196 ( .A0(conv_1[503]), .A1(n23430), .B0(n34666), .C0(n23429), 
        .Y(n23431) );
  OAI211XL U28197 ( .A0(n33427), .A1(n23432), .B0(n16652), .C0(n23431), .Y(
        n15960) );
  NAND2XL U28198 ( .A(n24217), .B(conv_1[195]), .Y(n24216) );
  INVXL U28199 ( .A(n24216), .Y(n23433) );
  NAND2XL U28200 ( .A(n23433), .B(n27429), .Y(n23434) );
  NAND2XL U28201 ( .A(n24221), .B(conv_1[196]), .Y(n24220) );
  NAND2XL U28202 ( .A(n23434), .B(n24220), .Y(n24141) );
  AOI222XL U28203 ( .A0(n24142), .A1(conv_1[197]), .B0(n24142), .B1(n24141), 
        .C0(conv_1[197]), .C1(n24141), .Y(n23436) );
  NAND2XL U28204 ( .A(n27231), .B(n27849), .Y(n23435) );
  NAND2XL U28205 ( .A(conv_1[200]), .B(n23441), .Y(n23440) );
  OAI211XL U28206 ( .A0(conv_1[200]), .A1(n23441), .B0(n33822), .C0(n23440), 
        .Y(n23442) );
  OAI211XL U28207 ( .A0(n35384), .A1(n23443), .B0(n34544), .C0(n23442), .Y(
        n16263) );
  NAND2XL U28208 ( .A(conv_1[201]), .B(n23682), .Y(n23449) );
  AOI21XL U28209 ( .A0(n34060), .A1(n23449), .B0(n23451), .Y(n23447) );
  NAND2XL U28210 ( .A(conv_1[202]), .B(n23447), .Y(n23446) );
  OAI211XL U28211 ( .A0(conv_1[202]), .A1(n23447), .B0(n33788), .C0(n23446), 
        .Y(n23448) );
  OAI211XL U28212 ( .A0(n35384), .A1(n23450), .B0(n16652), .C0(n23448), .Y(
        n16261) );
  NAND2XL U28213 ( .A(conv_1[203]), .B(n35372), .Y(n31111) );
  AOI21XL U28214 ( .A0(n34060), .A1(n31111), .B0(n31113), .Y(n23453) );
  NAND2XL U28215 ( .A(conv_1[204]), .B(n23453), .Y(n23452) );
  OAI211XL U28216 ( .A0(conv_1[204]), .A1(n23453), .B0(n16657), .C0(n23452), 
        .Y(n23454) );
  OAI211XL U28217 ( .A0(n35384), .A1(n31112), .B0(n16652), .C0(n23454), .Y(
        n16259) );
  OAI2BB1XL U28218 ( .A0N(n23457), .A1N(n23459), .B0(n23456), .Y(n23458) );
  OAI211XL U28219 ( .A0(n35986), .A1(n23459), .B0(n23458), .C0(n35847), .Y(
        n15326) );
  OR2XL U28220 ( .A(n23460), .B(n28721), .Y(n33524) );
  INVXL U28221 ( .A(n23463), .Y(n23465) );
  NAND2XL U28222 ( .A(n33403), .B(n23465), .Y(n23464) );
  OAI31XL U28223 ( .A0(n33403), .A1(n28721), .A2(n23465), .B0(n23464), .Y(
        n23966) );
  NAND2XL U28224 ( .A(n23966), .B(conv_1[257]), .Y(n23965) );
  NAND2BXL U28225 ( .AN(n23466), .B(n23965), .Y(n23468) );
  NOR2X1 U28226 ( .A(n23467), .B(n23468), .Y(n24688) );
  NAND2XL U28227 ( .A(conv_1[258]), .B(n23470), .Y(n23469) );
  OAI211XL U28228 ( .A0(conv_1[258]), .A1(n23470), .B0(n16656), .C0(n23469), 
        .Y(n23471) );
  OAI211XL U28229 ( .A0(n34080), .A1(n23472), .B0(n32867), .C0(n23471), .Y(
        n16205) );
  INVXL U28230 ( .A(conv_2[79]), .Y(n23484) );
  NAND2XL U28231 ( .A(n29046), .B(n34438), .Y(n23480) );
  INVXL U28232 ( .A(conv_2[75]), .Y(n34439) );
  NAND2XL U28233 ( .A(n23473), .B(n34436), .Y(n23475) );
  INVXL U28234 ( .A(n34436), .Y(n23474) );
  AOI221XL U28235 ( .A0(n18913), .A1(n23474), .B0(n28126), .B1(n34436), .C0(
        n33020), .Y(n23947) );
  NAND2XL U28236 ( .A(n23947), .B(conv_2[76]), .Y(n23946) );
  NAND2XL U28237 ( .A(n28128), .B(n23477), .Y(n23478) );
  NAND2XL U28238 ( .A(n35853), .B(n23477), .Y(n23476) );
  NAND2XL U28239 ( .A(n30418), .B(conv_2[77]), .Y(n30417) );
  NAND2XL U28240 ( .A(conv_2[79]), .B(n23482), .Y(n23481) );
  OAI211XL U28241 ( .A0(conv_2[79]), .A1(n23482), .B0(n31735), .C0(n23481), 
        .Y(n23483) );
  OAI211XL U28242 ( .A0(n35879), .A1(n23484), .B0(n34408), .C0(n23483), .Y(
        n15234) );
  INVXL U28243 ( .A(conv_3[303]), .Y(n23490) );
  XOR2XL U28244 ( .A(n23486), .B(n23485), .Y(n23488) );
  NAND2XL U28245 ( .A(conv_3[303]), .B(n23488), .Y(n23487) );
  OAI211XL U28246 ( .A0(conv_3[303]), .A1(n23488), .B0(n31735), .C0(n23487), 
        .Y(n23489) );
  OAI211XL U28247 ( .A0(n35736), .A1(n23490), .B0(n35574), .C0(n23489), .Y(
        n15795) );
  INVXL U28248 ( .A(conv_3[273]), .Y(n23497) );
  AOI21XL U28249 ( .A0(n23493), .A1(n23492), .B0(n23491), .Y(n23495) );
  NAND2XL U28250 ( .A(conv_3[273]), .B(n23495), .Y(n23494) );
  OAI211XL U28251 ( .A0(conv_3[273]), .A1(n23495), .B0(n31735), .C0(n23494), 
        .Y(n23496) );
  OAI211XL U28252 ( .A0(n34709), .A1(n23497), .B0(n35574), .C0(n23496), .Y(
        n15797) );
  INVXL U28253 ( .A(conv_3[363]), .Y(n23503) );
  NOR2X1 U28254 ( .A(n27620), .B(n23504), .Y(n31330) );
  OAI21XL U28255 ( .A0(n30536), .A1(n23504), .B0(n31329), .Y(n23498) );
  INVXL U28256 ( .A(n23498), .Y(n30563) );
  AOI21XL U28257 ( .A0(n23505), .A1(n23506), .B0(n23499), .Y(n23501) );
  NAND2XL U28258 ( .A(conv_3[363]), .B(n23501), .Y(n23500) );
  OAI211XL U28259 ( .A0(conv_3[363]), .A1(n23501), .B0(n31735), .C0(n23500), 
        .Y(n23502) );
  OAI211XL U28260 ( .A0(n35764), .A1(n23503), .B0(n35574), .C0(n23502), .Y(
        n15791) );
  INVXL U28261 ( .A(conv_3[364]), .Y(n23513) );
  AOI222XL U28262 ( .A0(n23506), .A1(n23505), .B0(n23506), .B1(conv_3[363]), 
        .C0(n23505), .C1(conv_3[363]), .Y(n23507) );
  INVXL U28263 ( .A(n23507), .Y(n23508) );
  NAND2XL U28264 ( .A(conv_3[364]), .B(n23511), .Y(n23510) );
  OAI211XL U28265 ( .A0(conv_3[364]), .A1(n23511), .B0(n32611), .C0(n23510), 
        .Y(n23512) );
  OAI211XL U28266 ( .A0(n35764), .A1(n23513), .B0(n34097), .C0(n23512), .Y(
        n15755) );
  INVXL U28267 ( .A(conv_3[484]), .Y(n23521) );
  AND2XL U28268 ( .A(n23517), .B(n23516), .Y(n23773) );
  NAND2XL U28269 ( .A(conv_3[484]), .B(n23519), .Y(n23518) );
  OAI211XL U28270 ( .A0(conv_3[484]), .A1(n23519), .B0(n36020), .C0(n23518), 
        .Y(n23520) );
  OAI211XL U28271 ( .A0(n35826), .A1(n23521), .B0(n23520), .C0(n34097), .Y(
        n15747) );
  INVXL U28272 ( .A(conv_3[138]), .Y(n23530) );
  NAND4XL U28273 ( .A(conv_3[135]), .B(n29680), .C(n29678), .D(n34740), .Y(
        n23523) );
  NAND2XL U28274 ( .A(conv_3[135]), .B(n29678), .Y(n23522) );
  INVXL U28275 ( .A(n23522), .Y(n34738) );
  AOI221XL U28276 ( .A0(n30536), .A1(n23522), .B0(n29680), .B1(n34738), .C0(
        n34426), .Y(n27524) );
  NAND2XL U28277 ( .A(n27524), .B(conv_3[136]), .Y(n27523) );
  NAND2XL U28278 ( .A(n23523), .B(n27523), .Y(n23524) );
  NAND2XL U28279 ( .A(n27619), .B(n23524), .Y(n30708) );
  AOI2BB1XL U28280 ( .A0N(n18997), .A1N(n34426), .B0(n23524), .Y(n23525) );
  INVXL U28281 ( .A(n23525), .Y(n30707) );
  NAND2XL U28282 ( .A(conv_3[137]), .B(n30707), .Y(n23526) );
  NAND2XL U28283 ( .A(n30708), .B(n23526), .Y(n23531) );
  XOR2XL U28284 ( .A(n23532), .B(n23531), .Y(n23528) );
  NAND2XL U28285 ( .A(conv_3[138]), .B(n23528), .Y(n23527) );
  OAI211XL U28286 ( .A0(conv_3[138]), .A1(n23528), .B0(n32052), .C0(n23527), 
        .Y(n23529) );
  OAI211XL U28287 ( .A0(n34737), .A1(n23530), .B0(n35574), .C0(n23529), .Y(
        n15806) );
  INVXL U28288 ( .A(conv_3[139]), .Y(n23538) );
  NAND2XL U28289 ( .A(n24467), .B(n34740), .Y(n23534) );
  AOI222XL U28290 ( .A0(n23532), .A1(conv_3[138]), .B0(n23532), .B1(n23531), 
        .C0(conv_3[138]), .C1(n23531), .Y(n23533) );
  NAND2XL U28291 ( .A(n23534), .B(n23533), .Y(n23776) );
  NOR2BXL U28292 ( .AN(n23776), .B(n23777), .Y(n23536) );
  NAND2XL U28293 ( .A(conv_3[139]), .B(n23536), .Y(n23535) );
  OAI211XL U28294 ( .A0(conv_3[139]), .A1(n23536), .B0(n35336), .C0(n23535), 
        .Y(n23537) );
  OAI211XL U28295 ( .A0(n34737), .A1(n23538), .B0(n34097), .C0(n23537), .Y(
        n15770) );
  INVXL U28296 ( .A(conv_1[198]), .Y(n23544) );
  NAND2XL U28297 ( .A(conv_1[198]), .B(n23542), .Y(n23541) );
  OAI211XL U28298 ( .A0(conv_1[198]), .A1(n23542), .B0(n24499), .C0(n23541), 
        .Y(n23543) );
  OAI211XL U28299 ( .A0(n35384), .A1(n23544), .B0(n32867), .C0(n23543), .Y(
        n16265) );
  INVXL U28300 ( .A(conv_3[539]), .Y(n31290) );
  INVXL U28301 ( .A(conv_3[529]), .Y(n23554) );
  NAND2XL U28302 ( .A(conv_3[525]), .B(n29678), .Y(n23545) );
  NAND2XL U28303 ( .A(n28620), .B(n29680), .Y(n33328) );
  AOI21XL U28304 ( .A0(n30536), .A1(n23545), .B0(n33429), .Y(n33329) );
  NAND2XL U28305 ( .A(conv_3[526]), .B(n33329), .Y(n33326) );
  NAND2XL U28306 ( .A(n33328), .B(n33326), .Y(n23547) );
  NAND2XL U28307 ( .A(n18997), .B(n23547), .Y(n23546) );
  OAI31XL U28308 ( .A0(n18997), .A1(n33429), .A2(n23547), .B0(n23546), .Y(
        n30504) );
  NAND2XL U28309 ( .A(n23547), .B(n27619), .Y(n23548) );
  OAI2BB1XL U28310 ( .A0N(conv_3[527]), .A1N(n30504), .B0(n23548), .Y(n23734)
         );
  AND2XL U28311 ( .A(n23550), .B(n23549), .Y(n24365) );
  NAND2XL U28312 ( .A(conv_3[529]), .B(n23552), .Y(n23551) );
  OAI211XL U28313 ( .A0(conv_3[529]), .A1(n23552), .B0(n35336), .C0(n23551), 
        .Y(n23553) );
  OAI211XL U28314 ( .A0(n31191), .A1(n23554), .B0(n23553), .C0(n34097), .Y(
        n15744) );
  NAND2XL U28315 ( .A(conv_3[240]), .B(n30603), .Y(n30602) );
  INVXL U28316 ( .A(n33547), .Y(n33549) );
  OAI21XL U28317 ( .A0(n30536), .A1(n24021), .B0(n30602), .Y(n33548) );
  NAND2XL U28318 ( .A(conv_3[241]), .B(n33548), .Y(n33546) );
  NAND2XL U28319 ( .A(n33549), .B(n33546), .Y(n24022) );
  AOI22XL U28320 ( .A0(n32660), .A1(n23555), .B0(conv_3[242]), .B1(n33545), 
        .Y(n23556) );
  NAND2XL U28321 ( .A(n23556), .B(n35566), .Y(n15835) );
  ADDFXL U28322 ( .A(conv_3[182]), .B(n23558), .CI(n23557), .CO(n29733), .S(
        n23559) );
  AOI22XL U28323 ( .A0(n32660), .A1(n23559), .B0(conv_3[182]), .B1(n32650), 
        .Y(n23560) );
  NAND2XL U28324 ( .A(n23560), .B(n35566), .Y(n15839) );
  AOI22XL U28325 ( .A0(n33788), .A1(n23563), .B0(conv_3[362]), .B1(n33828), 
        .Y(n23564) );
  NAND2XL U28326 ( .A(n23564), .B(n35566), .Y(n15827) );
  OAI21XL U28327 ( .A0(n18913), .A1(n27764), .B0(n23565), .Y(n29800) );
  OR2XL U28328 ( .A(n23565), .B(n18913), .Y(n29799) );
  OAI2BB1XL U28329 ( .A0N(conv_2[511]), .A1N(n29800), .B0(n29799), .Y(n27765)
         );
  AOI22XL U28330 ( .A0(n32660), .A1(n23566), .B0(conv_2[512]), .B1(n33575), 
        .Y(n23567) );
  NAND2XL U28331 ( .A(n23567), .B(n34621), .Y(n15277) );
  NAND2XL U28332 ( .A(conv_2[180]), .B(n28124), .Y(n23568) );
  AOI221XL U28333 ( .A0(n34510), .A1(n28126), .B0(n23568), .B1(n18913), .C0(
        n34703), .Y(n31057) );
  NAND2XL U28334 ( .A(n34510), .B(n28126), .Y(n23569) );
  OAI2BB1XL U28335 ( .A0N(conv_2[181]), .A1N(n31057), .B0(n23569), .Y(n27081)
         );
  AOI22XL U28336 ( .A0(n33712), .A1(n23570), .B0(conv_2[182]), .B1(n33453), 
        .Y(n23571) );
  NAND2XL U28337 ( .A(n23571), .B(n34621), .Y(n15299) );
  NOR2X1 U28338 ( .A(n35853), .B(n34715), .Y(n25676) );
  OAI22XL U28339 ( .A0(n18913), .A1(n23574), .B0(n23573), .B1(n23572), .Y(
        n25675) );
  AOI22XL U28340 ( .A0(n33712), .A1(n23576), .B0(conv_2[107]), .B1(n23575), 
        .Y(n23577) );
  NAND2XL U28341 ( .A(n23577), .B(n34621), .Y(n15304) );
  INVXL U28342 ( .A(conv_2[29]), .Y(n27942) );
  NAND2XL U28343 ( .A(n34721), .B(n28068), .Y(n23581) );
  NAND2XL U28344 ( .A(n24199), .B(conv_2[15]), .Y(n24198) );
  INVXL U28345 ( .A(n24198), .Y(n23578) );
  NAND2XL U28346 ( .A(n23578), .B(n28126), .Y(n23579) );
  OAI32XL U28347 ( .A0(n18913), .A1(n30195), .A2(n23578), .B0(n24198), .B1(
        n28126), .Y(n24213) );
  NAND2XL U28348 ( .A(n24213), .B(conv_2[16]), .Y(n24212) );
  AOI222XL U28349 ( .A0(n30407), .A1(conv_2[17]), .B0(n30407), .B1(n30406), 
        .C0(conv_2[17]), .C1(n30406), .Y(n23580) );
  NAND2XL U28350 ( .A(conv_2[18]), .B(n23583), .Y(n23582) );
  OAI211XL U28351 ( .A0(conv_2[18]), .A1(n23583), .B0(n16657), .C0(n23582), 
        .Y(n23584) );
  OAI211XL U28352 ( .A0(n30412), .A1(n23585), .B0(n34105), .C0(n23584), .Y(
        n15274) );
  NAND2XL U28353 ( .A(n27231), .B(n34706), .Y(n23589) );
  OR2XL U28354 ( .A(n24137), .B(n35272), .Y(n23587) );
  NAND2XL U28355 ( .A(n24137), .B(n27429), .Y(n23586) );
  NAND2XL U28356 ( .A(n24148), .B(conv_1[181]), .Y(n24147) );
  AOI222XL U28357 ( .A0(n23970), .A1(conv_1[182]), .B0(n23970), .B1(n23969), 
        .C0(conv_1[182]), .C1(n23969), .Y(n23588) );
  NAND2XL U28358 ( .A(conv_1[186]), .B(n35352), .Y(n23597) );
  AOI21XL U28359 ( .A0(n32988), .A1(n23597), .B0(n23599), .Y(n23595) );
  NAND2XL U28360 ( .A(conv_1[187]), .B(n23595), .Y(n23594) );
  OAI211XL U28361 ( .A0(conv_1[187]), .A1(n23595), .B0(n33778), .C0(n23594), 
        .Y(n23596) );
  OAI211XL U28362 ( .A0(n35368), .A1(n23598), .B0(n34544), .C0(n23596), .Y(
        n16276) );
  NAND2XL U28363 ( .A(conv_1[188]), .B(n35358), .Y(n25063) );
  AOI21XL U28364 ( .A0(n32988), .A1(n25063), .B0(n25062), .Y(n23601) );
  NAND2XL U28365 ( .A(conv_1[189]), .B(n23601), .Y(n23600) );
  OAI211XL U28366 ( .A0(conv_1[189]), .A1(n23601), .B0(n33778), .C0(n23600), 
        .Y(n23602) );
  OAI211XL U28367 ( .A0(n35368), .A1(n25064), .B0(n16652), .C0(n23602), .Y(
        n16274) );
  INVXL U28368 ( .A(conv_3[333]), .Y(n23610) );
  NAND2XL U28369 ( .A(n29677), .B(n34525), .Y(n23606) );
  NAND2XL U28370 ( .A(n30615), .B(conv_3[330]), .Y(n30614) );
  INVXL U28371 ( .A(n30614), .Y(n23603) );
  NAND2XL U28372 ( .A(n23603), .B(n29680), .Y(n23604) );
  OAI32XL U28373 ( .A0(n23603), .A1(n34522), .A2(n30536), .B0(n29680), .B1(
        n30614), .Y(n30599) );
  NAND2XL U28374 ( .A(n30599), .B(conv_3[331]), .Y(n30598) );
  AOI222XL U28375 ( .A0(n30623), .A1(conv_3[332]), .B0(n30623), .B1(n30622), 
        .C0(conv_3[332]), .C1(n30622), .Y(n23605) );
  NAND2XL U28376 ( .A(n23606), .B(n23605), .Y(n23765) );
  NOR2BXL U28377 ( .AN(n23765), .B(n23766), .Y(n23608) );
  NAND2XL U28378 ( .A(conv_3[333]), .B(n23608), .Y(n23607) );
  OAI211XL U28379 ( .A0(conv_3[333]), .A1(n23608), .B0(n31735), .C0(n23607), 
        .Y(n23609) );
  OAI211XL U28380 ( .A0(n35748), .A1(n23610), .B0(n23609), .C0(n35574), .Y(
        n15793) );
  INVXL U28381 ( .A(conv_1[183]), .Y(n23616) );
  NAND2XL U28382 ( .A(conv_1[183]), .B(n23614), .Y(n23613) );
  OAI211XL U28383 ( .A0(conv_1[183]), .A1(n23614), .B0(n33778), .C0(n23613), 
        .Y(n23615) );
  OAI211XL U28384 ( .A0(n35368), .A1(n23616), .B0(n32867), .C0(n23615), .Y(
        n16280) );
  NAND2XL U28385 ( .A(conv_3[210]), .B(n29678), .Y(n23617) );
  NAND2XL U28386 ( .A(n27492), .B(n29680), .Y(n30530) );
  AOI21XL U28387 ( .A0(n30536), .A1(n23617), .B0(n28660), .Y(n30531) );
  NAND2XL U28388 ( .A(conv_3[211]), .B(n30531), .Y(n23618) );
  NAND2XL U28389 ( .A(n30530), .B(n23618), .Y(n23620) );
  NAND2XL U28390 ( .A(n18997), .B(n23620), .Y(n23619) );
  OAI31XL U28391 ( .A0(n18997), .A1(n28660), .A2(n23620), .B0(n23619), .Y(
        n30629) );
  NAND2XL U28392 ( .A(n23620), .B(n27619), .Y(n23621) );
  OAI2BB1XL U28393 ( .A0N(conv_3[212]), .A1N(n30629), .B0(n23621), .Y(n24322)
         );
  NAND2XL U28394 ( .A(conv_3[214]), .B(n23625), .Y(n23624) );
  OAI211XL U28395 ( .A0(conv_3[214]), .A1(n23625), .B0(n35336), .C0(n23624), 
        .Y(n23626) );
  OAI211XL U28396 ( .A0(n35665), .A1(n23627), .B0(n34097), .C0(n23626), .Y(
        n15765) );
  INVXL U28397 ( .A(conv_3[404]), .Y(n34009) );
  INVXL U28398 ( .A(conv_3[394]), .Y(n23637) );
  NAND4XL U28399 ( .A(conv_3[390]), .B(n29680), .C(n29678), .D(n27990), .Y(
        n23629) );
  NAND2XL U28400 ( .A(conv_3[390]), .B(n29678), .Y(n23628) );
  INVXL U28401 ( .A(n23628), .Y(n27988) );
  AOI221XL U28402 ( .A0(n30536), .A1(n23628), .B0(n29680), .B1(n27988), .C0(
        n32016), .Y(n31035) );
  NAND2XL U28403 ( .A(n31035), .B(conv_3[391]), .Y(n31034) );
  NAND2XL U28404 ( .A(n23629), .B(n31034), .Y(n30851) );
  AOI222XL U28405 ( .A0(n30852), .A1(conv_3[392]), .B0(n30852), .B1(n30851), 
        .C0(conv_3[392]), .C1(n30851), .Y(n23631) );
  NAND2XL U28406 ( .A(n29677), .B(n27990), .Y(n23630) );
  NAND2XL U28407 ( .A(conv_3[394]), .B(n23635), .Y(n23634) );
  OAI211XL U28408 ( .A0(conv_3[394]), .A1(n23635), .B0(n35336), .C0(n23634), 
        .Y(n23636) );
  OAI211XL U28409 ( .A0(n33703), .A1(n23637), .B0(n34097), .C0(n23636), .Y(
        n15753) );
  NAND2XL U28410 ( .A(n27231), .B(n34224), .Y(n23640) );
  NAND2XL U28411 ( .A(n30663), .B(conv_1[435]), .Y(n30662) );
  OR2XL U28412 ( .A(n30662), .B(n35272), .Y(n30657) );
  OAI21XL U28413 ( .A0(n35272), .A1(n27898), .B0(n30662), .Y(n30656) );
  NAND2XL U28414 ( .A(conv_1[436]), .B(n30656), .Y(n23638) );
  NAND2XL U28415 ( .A(n30657), .B(n23638), .Y(n30580) );
  AOI222XL U28416 ( .A0(n30581), .A1(conv_1[437]), .B0(n30581), .B1(n30580), 
        .C0(conv_1[437]), .C1(n30580), .Y(n23639) );
  AND2XL U28417 ( .A(n23640), .B(n23639), .Y(n26940) );
  INVXL U28418 ( .A(n35515), .Y(n27149) );
  OAI21XL U28419 ( .A0(conv_1[441]), .A1(n27154), .B0(n35515), .Y(n25231) );
  INVXL U28420 ( .A(conv_1[442]), .Y(n25236) );
  INVXL U28421 ( .A(conv_1[440]), .Y(n27171) );
  AOI21XL U28422 ( .A0(n27155), .A1(conv_1[441]), .B0(n35515), .Y(n25232) );
  AOI22XL U28423 ( .A0(n24378), .A1(n23644), .B0(conv_1[443]), .B1(n35517), 
        .Y(n23645) );
  NAND2XL U28424 ( .A(n23645), .B(n34689), .Y(n16020) );
  ADDFX1 U28425 ( .A(conv_1[123]), .B(n23647), .CI(n23646), .CO(n23648), .S(
        n22431) );
  NOR2X1 U28426 ( .A(n23649), .B(n23648), .Y(n30754) );
  OAI31XL U28427 ( .A0(conv_1[127]), .A1(conv_1[128]), .A2(n34289), .B0(n34292), .Y(n26709) );
  NOR2X1 U28428 ( .A(n34292), .B(n34289), .Y(n29390) );
  INVXL U28429 ( .A(conv_1[127]), .Y(n29394) );
  AOI21XL U28430 ( .A0(conv_1[128]), .A1(n34291), .B0(n34292), .Y(n26710) );
  AOI22XL U28431 ( .A0(n32656), .A1(n23651), .B0(conv_1[130]), .B1(n23883), 
        .Y(n23652) );
  NAND2XL U28432 ( .A(n23652), .B(n34696), .Y(n16333) );
  ADDFXL U28433 ( .A(conv_1[502]), .B(n27131), .CI(n23653), .CO(n27119), .S(
        n23654) );
  AOI22XL U28434 ( .A0(n24378), .A1(n23654), .B0(conv_1[502]), .B1(n23663), 
        .Y(n23655) );
  NAND2XL U28435 ( .A(n23655), .B(n34544), .Y(n15961) );
  ADDFXL U28436 ( .A(conv_1[126]), .B(n34292), .CI(n23656), .CO(n34289), .S(
        n23657) );
  AOI22XL U28437 ( .A0(n32656), .A1(n23657), .B0(conv_1[126]), .B1(n23883), 
        .Y(n23658) );
  NAND2XL U28438 ( .A(n23658), .B(n34696), .Y(n16337) );
  AOI22XL U28439 ( .A0(n32656), .A1(n23660), .B0(conv_1[248]), .B1(n33658), 
        .Y(n23661) );
  NAND2XL U28440 ( .A(n23661), .B(n34682), .Y(n16215) );
  ADDFXL U28441 ( .A(conv_1[500]), .B(n27131), .CI(n23662), .CO(n26335), .S(
        n23664) );
  AOI22XL U28442 ( .A0(n24378), .A1(n23664), .B0(conv_1[500]), .B1(n23663), 
        .Y(n23665) );
  NAND2XL U28443 ( .A(n23665), .B(n34544), .Y(n15963) );
  INVXL U28444 ( .A(conv_3[288]), .Y(n23671) );
  NAND2XL U28445 ( .A(conv_3[288]), .B(n23669), .Y(n23668) );
  OAI211XL U28446 ( .A0(conv_3[288]), .A1(n23669), .B0(n31735), .C0(n23668), 
        .Y(n23670) );
  OAI211XL U28447 ( .A0(n35726), .A1(n23671), .B0(n35574), .C0(n23670), .Y(
        n15796) );
  AOI22XL U28448 ( .A0(n22896), .A1(n23674), .B0(n23673), .B1(n23672), .Y(
        N17505) );
  INVXL U28449 ( .A(conv_1[331]), .Y(n23678) );
  NAND2XL U28450 ( .A(conv_1[331]), .B(n23676), .Y(n23675) );
  OAI211XL U28451 ( .A0(conv_1[331]), .A1(n23676), .B0(n27932), .C0(n23675), 
        .Y(n23677) );
  OAI211XL U28452 ( .A0(n35437), .A1(n23678), .B0(n23677), .C0(n33067), .Y(
        n16132) );
  AOI221XL U28453 ( .A0(n23680), .A1(n33982), .B0(n23679), .B1(n16657), .C0(
        n35374), .Y(n23685) );
  OAI211XL U28454 ( .A0(n35379), .A1(n23682), .B0(n32611), .C0(n23681), .Y(
        n23683) );
  OAI211XL U28455 ( .A0(n23685), .A1(n23684), .B0(n16652), .C0(n23683), .Y(
        n16262) );
  INVXL U28456 ( .A(conv_3[134]), .Y(n34788) );
  INVXL U28457 ( .A(conv_3[124]), .Y(n23694) );
  OAI21XL U28458 ( .A0(n30536), .A1(n28948), .B0(n30837), .Y(n27514) );
  OAI21XL U28459 ( .A0(n18997), .A1(n28948), .B0(n23686), .Y(n23687) );
  INVXL U28460 ( .A(n23687), .Y(n30742) );
  INVXL U28461 ( .A(n23688), .Y(n23689) );
  NAND2XL U28462 ( .A(conv_3[124]), .B(n23692), .Y(n23691) );
  OAI211XL U28463 ( .A0(conv_3[124]), .A1(n23692), .B0(n35336), .C0(n23691), 
        .Y(n23693) );
  OAI211XL U28464 ( .A0(n35626), .A1(n23694), .B0(n34097), .C0(n23693), .Y(
        n15771) );
  AOI22XL U28465 ( .A0(n24378), .A1(intadd_2_SUM_1_), .B0(conv_1[3]), .B1(
        n24536), .Y(n23695) );
  NAND2XL U28466 ( .A(n23695), .B(n32867), .Y(n16460) );
  INVXL U28467 ( .A(conv_1[530]), .Y(n23700) );
  AOI211XL U28468 ( .A0(n23700), .A1(n23698), .B0(n36042), .C0(n23697), .Y(
        n23699) );
  AOI2BB1XL U28469 ( .A0N(n23700), .A1N(n33432), .B0(n23699), .Y(n23701) );
  NAND2XL U28470 ( .A(n23701), .B(n34682), .Y(n15933) );
  ADDFXL U28471 ( .A(conv_2[273]), .B(n23703), .CI(n23702), .CO(n29063), .S(
        n23704) );
  AOI22XL U28472 ( .A0(n24378), .A1(n23704), .B0(conv_2[273]), .B1(n35952), 
        .Y(n23705) );
  NAND2XL U28473 ( .A(n23705), .B(n34105), .Y(n15257) );
  NAND2XL U28474 ( .A(conv_2[210]), .B(n28124), .Y(n23706) );
  AOI21XL U28475 ( .A0(n18913), .A1(n23706), .B0(n28660), .Y(n31047) );
  NAND2XL U28476 ( .A(n34473), .B(n28126), .Y(n31046) );
  OAI2BB1XL U28477 ( .A0N(conv_2[211]), .A1N(n31047), .B0(n31046), .Y(n23708)
         );
  NAND2XL U28478 ( .A(n35853), .B(n23708), .Y(n23707) );
  NAND2XL U28479 ( .A(n23708), .B(n28128), .Y(n23709) );
  OAI2BB1XL U28480 ( .A0N(conv_2[212]), .A1N(n27051), .B0(n23709), .Y(n28661)
         );
  AOI22XL U28481 ( .A0(n24378), .A1(n23710), .B0(conv_2[213]), .B1(n33765), 
        .Y(n23711) );
  NAND2XL U28482 ( .A(n23711), .B(n34105), .Y(n15261) );
  AOI22XL U28483 ( .A0(n24378), .A1(n23714), .B0(conv_2[348]), .B1(n24190), 
        .Y(n23715) );
  NAND2XL U28484 ( .A(n23715), .B(n34105), .Y(n15252) );
  NAND2XL U28485 ( .A(conv_2[450]), .B(n28124), .Y(n23716) );
  NAND2XL U28486 ( .A(n34442), .B(n28126), .Y(n29787) );
  AOI21XL U28487 ( .A0(n18913), .A1(n23716), .B0(n27644), .Y(n29788) );
  NAND2XL U28488 ( .A(conv_2[451]), .B(n29788), .Y(n23717) );
  NAND2XL U28489 ( .A(n29787), .B(n23717), .Y(n23719) );
  NAND2XL U28490 ( .A(n35853), .B(n23719), .Y(n23718) );
  NAND2XL U28491 ( .A(n23719), .B(n28128), .Y(n23720) );
  OAI2BB1XL U28492 ( .A0N(conv_2[452]), .A1N(n30015), .B0(n23720), .Y(n24337)
         );
  AOI22XL U28493 ( .A0(n24378), .A1(n23721), .B0(conv_2[453]), .B1(n33606), 
        .Y(n23722) );
  NAND2XL U28494 ( .A(n23722), .B(n34105), .Y(n15245) );
  INVXL U28495 ( .A(conv_1[377]), .Y(n23728) );
  NAND2XL U28496 ( .A(conv_1[377]), .B(n23726), .Y(n23725) );
  OAI211XL U28497 ( .A0(conv_1[377]), .A1(n23726), .B0(n34028), .C0(n23725), 
        .Y(n23727) );
  OAI211XL U28498 ( .A0(n35466), .A1(n23728), .B0(n33542), .C0(n23727), .Y(
        n16086) );
  ADDFXL U28499 ( .A(conv_3[78]), .B(n23730), .CI(n23729), .CO(n22920), .S(
        n23732) );
  AOI22XL U28500 ( .A0(n32656), .A1(n23732), .B0(conv_3[78]), .B1(n23731), .Y(
        n23733) );
  NAND2XL U28501 ( .A(n23733), .B(n35574), .Y(n15810) );
  AOI22XL U28502 ( .A0(n32611), .A1(n23736), .B0(conv_3[528]), .B1(n33714), 
        .Y(n23737) );
  NAND2XL U28503 ( .A(n23737), .B(n35574), .Y(n15780) );
  AOI22XL U28504 ( .A0(n32611), .A1(n23740), .B0(conv_3[513]), .B1(n24479), 
        .Y(n23741) );
  NAND2XL U28505 ( .A(n23741), .B(n35574), .Y(n15781) );
  OAI2BB1XL U28506 ( .A0N(n23746), .A1N(n23744), .B0(n23743), .Y(n23745) );
  OAI211XL U28507 ( .A0(n34392), .A1(n23746), .B0(n33550), .C0(n23745), .Y(
        n15884) );
  INVX1 U28508 ( .A(n22257), .Y(n34433) );
  NAND2XL U28509 ( .A(n29678), .B(conv_3[165]), .Y(n23747) );
  OR2XL U28510 ( .A(n23747), .B(n22257), .Y(n28762) );
  INVXL U28511 ( .A(conv_3[166]), .Y(n27483) );
  OAI2BB1XL U28512 ( .A0N(n30536), .A1N(n23747), .B0(n34433), .Y(n27479) );
  NOR2X1 U28513 ( .A(n27478), .B(n23748), .Y(n23749) );
  OAI2BB1XL U28514 ( .A0N(n27619), .A1N(n34433), .B0(n23749), .Y(n35557) );
  NOR2X1 U28515 ( .A(n18997), .B(n23749), .Y(n35554) );
  NOR2BXL U28516 ( .AN(n35557), .B(n35558), .Y(n29068) );
  AOI22XL U28517 ( .A0(n32611), .A1(n23750), .B0(conv_3[168]), .B1(n35641), 
        .Y(n23751) );
  NAND2XL U28518 ( .A(n23751), .B(n35574), .Y(n15804) );
  NAND2XL U28519 ( .A(n23752), .B(n29680), .Y(n23753) );
  OAI32XL U28520 ( .A0(n30536), .A1(n23752), .A2(n35857), .B0(n31026), .B1(
        n29680), .Y(n27510) );
  NAND2XL U28521 ( .A(conv_3[1]), .B(n27510), .Y(n27509) );
  NAND2XL U28522 ( .A(n18997), .B(n23755), .Y(n23754) );
  OAI31XL U28523 ( .A0(n18997), .A1(n35857), .A2(n23755), .B0(n23754), .Y(
        n30786) );
  NAND2XL U28524 ( .A(n23755), .B(n27619), .Y(n23756) );
  INVXL U28525 ( .A(conv_3[14]), .Y(n33160) );
  AOI22XL U28526 ( .A0(n32611), .A1(n23757), .B0(conv_3[4]), .B1(n27508), .Y(
        n23758) );
  NAND2XL U28527 ( .A(n23758), .B(n34097), .Y(n15779) );
  INVXL U28528 ( .A(conv_1[379]), .Y(n23764) );
  NAND2XL U28529 ( .A(conv_1[379]), .B(n23762), .Y(n23761) );
  OAI211XL U28530 ( .A0(conv_1[379]), .A1(n23762), .B0(n16657), .C0(n23761), 
        .Y(n23763) );
  OAI211XL U28531 ( .A0(n35466), .A1(n23764), .B0(n35489), .C0(n23763), .Y(
        n16084) );
  NAND2XL U28532 ( .A(n24467), .B(n34525), .Y(n23768) );
  NAND2XL U28533 ( .A(n23768), .B(n23767), .Y(n26946) );
  NAND2XL U28534 ( .A(n31967), .B(n23769), .Y(n35749) );
  AOI22XL U28535 ( .A0(n33712), .A1(n23770), .B0(conv_3[337]), .B1(n35756), 
        .Y(n23771) );
  NAND2XL U28536 ( .A(n23771), .B(n35588), .Y(n15521) );
  AOI22XL U28537 ( .A0(n33778), .A1(n23774), .B0(conv_3[485]), .B1(n35833), 
        .Y(n23775) );
  NAND2XL U28538 ( .A(n23775), .B(n35588), .Y(n15423) );
  NAND2XL U28539 ( .A(n32789), .B(n23778), .Y(n34396) );
  AOI21XL U28540 ( .A0(conv_3[140]), .A1(n34396), .B0(n33466), .Y(n31714) );
  AOI22XL U28541 ( .A0(n33778), .A1(n23779), .B0(conv_3[142]), .B1(n33461), 
        .Y(n23780) );
  NAND2XL U28542 ( .A(n23780), .B(n35588), .Y(n15651) );
  INVXL U28543 ( .A(conv_2[33]), .Y(n27704) );
  AOI22XL U28544 ( .A0(n23783), .A1(n23782), .B0(n34906), .B1(n23781), .Y(
        n23788) );
  NAND2XL U28545 ( .A(n33990), .B(n28126), .Y(n23790) );
  NAND2XL U28546 ( .A(conv_2[30]), .B(n28124), .Y(n33987) );
  NAND2XL U28547 ( .A(n18913), .B(n33987), .Y(n23791) );
  OAI211XL U28548 ( .A0(n18913), .A1(n33987), .B0(n33990), .C0(n23791), .Y(
        n24268) );
  INVXL U28549 ( .A(conv_2[31]), .Y(n24270) );
  OAI2BB1XL U28550 ( .A0N(n33990), .A1N(n28128), .B0(n23793), .Y(n31103) );
  AOI21XL U28551 ( .A0(conv_2[32]), .A1(n31103), .B0(n31102), .Y(n23795) );
  NAND2XL U28552 ( .A(n33990), .B(n28068), .Y(n23794) );
  AND2XL U28553 ( .A(n23795), .B(n23794), .Y(n27703) );
  NAND2XL U28554 ( .A(conv_2[33]), .B(n23797), .Y(n23796) );
  OAI211XL U28555 ( .A0(conv_2[33]), .A1(n23797), .B0(n33778), .C0(n23796), 
        .Y(n23798) );
  OAI211XL U28556 ( .A0(n35865), .A1(n27704), .B0(n34105), .C0(n23798), .Y(
        n15273) );
  INVXL U28557 ( .A(conv_2[480]), .Y(n23801) );
  OAI211XL U28558 ( .A0(n23799), .A1(conv_2[480]), .B0(n33982), .C0(n27734), 
        .Y(n23800) );
  OAI211XL U28559 ( .A0(n34137), .A1(n23801), .B0(n34583), .C0(n23800), .Y(
        n15351) );
  INVXL U28560 ( .A(conv_3[318]), .Y(n23809) );
  NAND2XL U28561 ( .A(n30611), .B(conv_3[315]), .Y(n30610) );
  OAI21XL U28562 ( .A0(n30536), .A1(n22269), .B0(n30610), .Y(n23802) );
  INVXL U28563 ( .A(n23802), .Y(n30557) );
  NAND2XL U28564 ( .A(n27619), .B(n23803), .Y(n35561) );
  INVXL U28565 ( .A(n35561), .Y(n35565) );
  INVXL U28566 ( .A(conv_3[317]), .Y(n35563) );
  NAND2XL U28567 ( .A(n23804), .B(n23805), .Y(n23810) );
  AND2XL U28568 ( .A(n23810), .B(n23811), .Y(n23807) );
  NAND2XL U28569 ( .A(conv_3[318]), .B(n23807), .Y(n23806) );
  OAI211XL U28570 ( .A0(conv_3[318]), .A1(n23807), .B0(n31735), .C0(n23806), 
        .Y(n23808) );
  OAI211XL U28571 ( .A0(n35743), .A1(n23809), .B0(n23808), .C0(n35574), .Y(
        n15794) );
  XOR2XL U28572 ( .A(n28756), .B(n28755), .Y(n23813) );
  NAND2XL U28573 ( .A(conv_3[319]), .B(n23813), .Y(n23812) );
  OAI211XL U28574 ( .A0(conv_3[319]), .A1(n23813), .B0(n32052), .C0(n23812), 
        .Y(n23814) );
  OAI211XL U28575 ( .A0(n35743), .A1(n23815), .B0(n23814), .C0(n34097), .Y(
        n15758) );
  INVXL U28576 ( .A(conv_1[375]), .Y(n23819) );
  OAI211XL U28577 ( .A0(n23817), .A1(conv_1[375]), .B0(n33982), .C0(n23816), 
        .Y(n23818) );
  OAI211XL U28578 ( .A0(n35466), .A1(n23819), .B0(n34773), .C0(n23818), .Y(
        n16088) );
  OAI2BB1XL U28579 ( .A0N(n23824), .A1N(n23822), .B0(n23821), .Y(n23823) );
  OAI211XL U28580 ( .A0(n35466), .A1(n23824), .B0(n33067), .C0(n23823), .Y(
        n16087) );
  INVXL U28581 ( .A(conv_2[46]), .Y(n23830) );
  NAND2XL U28582 ( .A(n23826), .B(n23825), .Y(n23828) );
  NAND2XL U28583 ( .A(n23830), .B(n23828), .Y(n23827) );
  OAI211XL U28584 ( .A0(n23830), .A1(n23828), .B0(n33982), .C0(n23827), .Y(
        n23829) );
  OAI211XL U28585 ( .A0(n34505), .A1(n23830), .B0(n23829), .C0(n35847), .Y(
        n15344) );
  INVXL U28586 ( .A(conv_2[60]), .Y(n23834) );
  OAI211XL U28587 ( .A0(conv_2[60]), .A1(n23832), .B0(n30090), .C0(n23831), 
        .Y(n23833) );
  OAI211XL U28588 ( .A0(n35846), .A1(n23834), .B0(n23833), .C0(n34583), .Y(
        n15379) );
  AOI21XL U28589 ( .A0(n35411), .A1(n33663), .B0(n23836), .Y(n23838) );
  NAND2XL U28590 ( .A(conv_1[249]), .B(n23838), .Y(n23837) );
  OAI211XL U28591 ( .A0(conv_1[249]), .A1(n23838), .B0(n33778), .C0(n23837), 
        .Y(n23839) );
  OAI211XL U28592 ( .A0(n35417), .A1(n23840), .B0(n34281), .C0(n23839), .Y(
        n16214) );
  NOR2BXL U28593 ( .AN(n23842), .B(n23841), .Y(n23844) );
  NAND2XL U28594 ( .A(conv_1[245]), .B(n23844), .Y(n23843) );
  OAI211XL U28595 ( .A0(conv_1[245]), .A1(n23844), .B0(n33778), .C0(n23843), 
        .Y(n23845) );
  OAI211XL U28596 ( .A0(n35417), .A1(n23846), .B0(n34696), .C0(n23845), .Y(
        n16218) );
  INVXL U28597 ( .A(conv_2[121]), .Y(n23852) );
  NAND2XL U28598 ( .A(n23848), .B(n23847), .Y(n23850) );
  NAND2XL U28599 ( .A(n23852), .B(n23850), .Y(n23849) );
  OAI211XL U28600 ( .A0(n23852), .A1(n23850), .B0(n30090), .C0(n23849), .Y(
        n23851) );
  OAI211XL U28601 ( .A0(n34491), .A1(n23852), .B0(n23851), .C0(n35847), .Y(
        n15339) );
  INVXL U28602 ( .A(conv_2[299]), .Y(n33300) );
  INVXL U28603 ( .A(conv_2[288]), .Y(n23861) );
  NAND4XL U28604 ( .A(conv_2[285]), .B(n28126), .C(n28124), .D(n34455), .Y(
        n23854) );
  NAND2XL U28605 ( .A(conv_2[285]), .B(n28124), .Y(n23853) );
  INVXL U28606 ( .A(n23853), .Y(n34453) );
  NAND2XL U28607 ( .A(n30303), .B(conv_2[286]), .Y(n30302) );
  NAND2XL U28608 ( .A(n23854), .B(n30302), .Y(n23856) );
  NAND2XL U28609 ( .A(n28128), .B(n23856), .Y(n23857) );
  NAND2XL U28610 ( .A(n35853), .B(n23856), .Y(n23855) );
  NAND2XL U28611 ( .A(n27412), .B(conv_2[287]), .Y(n27411) );
  XOR2XL U28612 ( .A(n28087), .B(n28086), .Y(n23859) );
  NAND2XL U28613 ( .A(conv_2[288]), .B(n23859), .Y(n23858) );
  OAI211XL U28614 ( .A0(conv_2[288]), .A1(n23859), .B0(n35336), .C0(n23858), 
        .Y(n23860) );
  OAI211XL U28615 ( .A0(n35963), .A1(n23861), .B0(n34105), .C0(n23860), .Y(
        n15256) );
  INVXL U28616 ( .A(conv_2[151]), .Y(n23865) );
  NAND2XL U28617 ( .A(conv_2[151]), .B(n23863), .Y(n23862) );
  OAI211XL U28618 ( .A0(conv_2[151]), .A1(n23863), .B0(n30090), .C0(n23862), 
        .Y(n23864) );
  OAI211XL U28619 ( .A0(n34631), .A1(n23865), .B0(n23864), .C0(n35847), .Y(
        n15337) );
  INVXL U28620 ( .A(conv_2[334]), .Y(n23872) );
  AOI21XL U28621 ( .A0(n23868), .A1(n23867), .B0(n23866), .Y(n23870) );
  NAND2XL U28622 ( .A(conv_2[334]), .B(n23870), .Y(n23869) );
  OAI211XL U28623 ( .A0(conv_2[334]), .A1(n23870), .B0(n33778), .C0(n23869), 
        .Y(n23871) );
  OAI211XL U28624 ( .A0(n36003), .A1(n23872), .B0(n34408), .C0(n23871), .Y(
        n15217) );
  NOR2BXL U28625 ( .AN(n23874), .B(n23873), .Y(n23876) );
  NAND2XL U28626 ( .A(conv_2[272]), .B(n23876), .Y(n23875) );
  OAI211XL U28627 ( .A0(conv_2[272]), .A1(n23876), .B0(n35336), .C0(n23875), 
        .Y(n23877) );
  OAI211XL U28628 ( .A0(n30994), .A1(n23878), .B0(n23877), .C0(n34621), .Y(
        n15293) );
  INVXL U28629 ( .A(conv_2[1]), .Y(n23882) );
  NAND2XL U28630 ( .A(conv_2[0]), .B(n24004), .Y(n35855) );
  INVXL U28631 ( .A(n35855), .Y(n23879) );
  OAI32XL U28632 ( .A0(n18913), .A1(n23879), .A2(n35857), .B0(n35855), .B1(
        n28126), .Y(n35854) );
  NAND2XL U28633 ( .A(conv_2[1]), .B(n35854), .Y(n23880) );
  OAI211XL U28634 ( .A0(conv_2[1]), .A1(n35854), .B0(n33982), .C0(n23880), .Y(
        n23881) );
  OAI211XL U28635 ( .A0(n30958), .A1(n23882), .B0(n23881), .C0(n35847), .Y(
        n15347) );
  OAI2BB1XL U28636 ( .A0N(n23886), .A1N(n23888), .B0(n23885), .Y(n23887) );
  OAI211XL U28637 ( .A0(n34296), .A1(n23888), .B0(n33067), .C0(n23887), .Y(
        n16342) );
  INVXL U28638 ( .A(conv_1[227]), .Y(n23894) );
  NAND2XL U28639 ( .A(n23890), .B(n23889), .Y(n23892) );
  NAND2XL U28640 ( .A(n23894), .B(n23892), .Y(n23891) );
  OAI211XL U28641 ( .A0(n23894), .A1(n23892), .B0(n24499), .C0(n23891), .Y(
        n23893) );
  OAI211XL U28642 ( .A0(n35408), .A1(n23894), .B0(n23893), .C0(n33542), .Y(
        n16236) );
  INVXL U28643 ( .A(conv_3[74]), .Y(n32168) );
  NAND2XL U28644 ( .A(n24467), .B(n34699), .Y(n23900) );
  NAND2XL U28645 ( .A(conv_3[60]), .B(n29678), .Y(n23895) );
  AOI221XL U28646 ( .A0(n34698), .A1(n29680), .B0(n23895), .B1(n30536), .C0(
        n31418), .Y(n27489) );
  NAND2XL U28647 ( .A(n34698), .B(n29680), .Y(n23896) );
  OAI2BB1XL U28648 ( .A0N(conv_3[61]), .A1N(n27489), .B0(n23896), .Y(n24236)
         );
  NAND2XL U28649 ( .A(n23898), .B(n23897), .Y(n34107) );
  OAI2BB1X1 U28650 ( .A0N(n34112), .A1N(n34107), .B0(n34108), .Y(n23899) );
  AND2X1 U28651 ( .A(n23900), .B(n23899), .Y(n31419) );
  NOR2X1 U28652 ( .A(n23900), .B(n23899), .Y(n31420) );
  NAND2XL U28653 ( .A(conv_3[64]), .B(n23902), .Y(n23901) );
  OAI211XL U28654 ( .A0(conv_3[64]), .A1(n23902), .B0(n35336), .C0(n23901), 
        .Y(n23903) );
  OAI211XL U28655 ( .A0(n35598), .A1(n23904), .B0(n34097), .C0(n23903), .Y(
        n15775) );
  INVXL U28656 ( .A(conv_1[212]), .Y(n23908) );
  NAND2XL U28657 ( .A(conv_1[212]), .B(n23906), .Y(n23905) );
  OAI211XL U28658 ( .A0(conv_1[212]), .A1(n23906), .B0(n16657), .C0(n23905), 
        .Y(n23907) );
  OAI211XL U28659 ( .A0(n35395), .A1(n23908), .B0(n23907), .C0(n33542), .Y(
        n16251) );
  NAND2XL U28660 ( .A(conv_1[229]), .B(n23912), .Y(n23911) );
  OAI211XL U28661 ( .A0(conv_1[229]), .A1(n23912), .B0(n33778), .C0(n23911), 
        .Y(n23913) );
  OAI211XL U28662 ( .A0(n35408), .A1(n23914), .B0(n23913), .C0(n35489), .Y(
        n16234) );
  INVXL U28663 ( .A(conv_1[177]), .Y(n23921) );
  AOI21XL U28664 ( .A0(n26667), .A1(n23923), .B0(n23917), .Y(n23919) );
  NAND2XL U28665 ( .A(conv_1[177]), .B(n23919), .Y(n23918) );
  OAI211XL U28666 ( .A0(conv_1[177]), .A1(n23919), .B0(n33778), .C0(n23918), 
        .Y(n23920) );
  OAI211XL U28667 ( .A0(n35346), .A1(n23921), .B0(n16652), .C0(n23920), .Y(
        n16286) );
  INVXL U28668 ( .A(conv_1[172]), .Y(n23927) );
  AOI21XL U28669 ( .A0(n27539), .A1(n23923), .B0(n23922), .Y(n23925) );
  NAND2XL U28670 ( .A(conv_1[172]), .B(n23925), .Y(n23924) );
  OAI211XL U28671 ( .A0(conv_1[172]), .A1(n23925), .B0(n24499), .C0(n23924), 
        .Y(n23926) );
  OAI211XL U28672 ( .A0(n35346), .A1(n23927), .B0(n34689), .C0(n23926), .Y(
        n16291) );
  INVXL U28673 ( .A(conv_3[50]), .Y(n34375) );
  OAI2BB1XL U28674 ( .A0N(conv_3[49]), .A1N(n23929), .B0(n23928), .Y(n23930)
         );
  NAND2XL U28675 ( .A(n33824), .B(n23930), .Y(n34371) );
  NAND2XL U28676 ( .A(n34375), .B(n34371), .Y(n31211) );
  OAI21XL U28677 ( .A0(conv_3[52]), .A1(n31204), .B0(n33824), .Y(n34387) );
  NAND2XL U28678 ( .A(n34393), .B(n34387), .Y(n23931) );
  OR2XL U28679 ( .A(n23930), .B(n33824), .Y(n34370) );
  AOI21XL U28680 ( .A0(conv_3[50]), .A1(n34370), .B0(n33824), .Y(n31210) );
  OAI2BB1XL U28681 ( .A0N(conv_3[52]), .A1N(n31205), .B0(n32178), .Y(n34386)
         );
  AND2XL U28682 ( .A(n23931), .B(n34386), .Y(n31199) );
  NAND2XL U28683 ( .A(n33824), .B(n23931), .Y(n31197) );
  OAI21XL U28684 ( .A0(n33824), .A1(n31199), .B0(n31197), .Y(n23933) );
  NAND2XL U28685 ( .A(n31198), .B(n23933), .Y(n23932) );
  OAI211XL U28686 ( .A0(n31198), .A1(n23933), .B0(n33778), .C0(n23932), .Y(
        n23934) );
  OAI211XL U28687 ( .A0(n34392), .A1(n31198), .B0(n35588), .C0(n23934), .Y(
        n15709) );
  INVXL U28688 ( .A(conv_1[174]), .Y(n23940) );
  NAND2XL U28689 ( .A(conv_1[174]), .B(n23938), .Y(n23937) );
  OAI211XL U28690 ( .A0(conv_1[174]), .A1(n23938), .B0(n33778), .C0(n23937), 
        .Y(n23939) );
  OAI211XL U28691 ( .A0(n35346), .A1(n23940), .B0(n16652), .C0(n23939), .Y(
        n16289) );
  OAI2BB1XL U28692 ( .A0N(n23945), .A1N(n23943), .B0(n23942), .Y(n23944) );
  OAI211XL U28693 ( .A0(n34271), .A1(n23945), .B0(n33067), .C0(n23944), .Y(
        n16327) );
  INVXL U28694 ( .A(conv_2[76]), .Y(n23949) );
  OAI211XL U28695 ( .A0(n23947), .A1(conv_2[76]), .B0(n33982), .C0(n23946), 
        .Y(n23948) );
  OAI211XL U28696 ( .A0(n35879), .A1(n23949), .B0(n35847), .C0(n23948), .Y(
        n15342) );
  OAI211XL U28697 ( .A0(n23951), .A1(conv_1[226]), .B0(n31735), .C0(n23950), 
        .Y(n23952) );
  OAI211XL U28698 ( .A0(n35408), .A1(n23953), .B0(n23952), .C0(n33067), .Y(
        n16237) );
  INVXL U28699 ( .A(conv_3[449]), .Y(n32149) );
  INVXL U28700 ( .A(conv_3[439]), .Y(n23964) );
  NAND2XL U28701 ( .A(n24467), .B(n34224), .Y(n23960) );
  NAND2XL U28702 ( .A(n29677), .B(n34224), .Y(n23958) );
  NAND2XL U28703 ( .A(n29678), .B(conv_3[435]), .Y(n23955) );
  INVXL U28704 ( .A(n23955), .Y(n34223) );
  NAND2XL U28705 ( .A(n23954), .B(n34223), .Y(n23956) );
  AOI221XL U28706 ( .A0(n30536), .A1(n23955), .B0(n29680), .B1(n34223), .C0(
        n27898), .Y(n31031) );
  NAND2XL U28707 ( .A(n31031), .B(conv_3[436]), .Y(n31030) );
  NAND2XL U28708 ( .A(n23956), .B(n31030), .Y(n30811) );
  AOI222XL U28709 ( .A0(n30812), .A1(conv_3[437]), .B0(n30812), .B1(n30811), 
        .C0(conv_3[437]), .C1(n30811), .Y(n23957) );
  NAND2XL U28710 ( .A(n23958), .B(n23957), .Y(n29708) );
  OAI21XL U28711 ( .A0(conv_3[438]), .A1(n29707), .B0(n29708), .Y(n23959) );
  NAND2XL U28712 ( .A(conv_3[439]), .B(n23962), .Y(n23961) );
  OAI211XL U28713 ( .A0(conv_3[439]), .A1(n23962), .B0(n36020), .C0(n23961), 
        .Y(n23963) );
  OAI211XL U28714 ( .A0(n35792), .A1(n23964), .B0(n34097), .C0(n23963), .Y(
        n15750) );
  OAI211XL U28715 ( .A0(n23966), .A1(conv_1[257]), .B0(n32660), .C0(n23965), 
        .Y(n23967) );
  OAI211XL U28716 ( .A0(n34080), .A1(n23968), .B0(n33542), .C0(n23967), .Y(
        n16206) );
  INVXL U28717 ( .A(conv_1[182]), .Y(n23974) );
  XOR2XL U28718 ( .A(n23970), .B(n23969), .Y(n23972) );
  NAND2XL U28719 ( .A(conv_1[182]), .B(n23972), .Y(n23971) );
  OAI211XL U28720 ( .A0(conv_1[182]), .A1(n23972), .B0(n33778), .C0(n23971), 
        .Y(n23973) );
  OAI211XL U28721 ( .A0(n35368), .A1(n23974), .B0(n33542), .C0(n23973), .Y(
        n16281) );
  INVXL U28722 ( .A(conv_1[184]), .Y(n23980) );
  NAND2XL U28723 ( .A(conv_1[184]), .B(n23978), .Y(n23977) );
  OAI211XL U28724 ( .A0(conv_1[184]), .A1(n23978), .B0(n33778), .C0(n23977), 
        .Y(n23979) );
  OAI211XL U28725 ( .A0(n35368), .A1(n23980), .B0(n35489), .C0(n23979), .Y(
        n16279) );
  INVXL U28726 ( .A(conv_1[316]), .Y(n23986) );
  NAND2XL U28727 ( .A(n23982), .B(n23981), .Y(n23984) );
  NAND2XL U28728 ( .A(n23986), .B(n23984), .Y(n23983) );
  OAI211XL U28729 ( .A0(n23986), .A1(n23984), .B0(n30090), .C0(n23983), .Y(
        n23985) );
  OAI211XL U28730 ( .A0(n34263), .A1(n23986), .B0(n23985), .C0(n33067), .Y(
        n16147) );
  INVXL U28731 ( .A(conv_2[375]), .Y(n23990) );
  OAI211XL U28732 ( .A0(n23988), .A1(conv_2[375]), .B0(n30090), .C0(n23987), 
        .Y(n23989) );
  OAI211XL U28733 ( .A0(n36028), .A1(n23990), .B0(n34583), .C0(n23989), .Y(
        n15358) );
  INVXL U28734 ( .A(conv_2[378]), .Y(n23996) );
  NAND2XL U28735 ( .A(conv_2[378]), .B(n23994), .Y(n23993) );
  OAI211XL U28736 ( .A0(conv_2[378]), .A1(n23994), .B0(n35336), .C0(n23993), 
        .Y(n23995) );
  OAI211XL U28737 ( .A0(n36028), .A1(n23996), .B0(n34105), .C0(n23995), .Y(
        n15250) );
  INVXL U28738 ( .A(conv_1[214]), .Y(n24003) );
  AOI21XL U28739 ( .A0(n23999), .A1(n23998), .B0(n23997), .Y(n24001) );
  NAND2XL U28740 ( .A(conv_1[214]), .B(n24001), .Y(n24000) );
  OAI211XL U28741 ( .A0(conv_1[214]), .A1(n24001), .B0(n33712), .C0(n24000), 
        .Y(n24002) );
  OAI211XL U28742 ( .A0(n35395), .A1(n24003), .B0(n35489), .C0(n24002), .Y(
        n16249) );
  OAI211XL U28743 ( .A0(conv_2[0]), .A1(n24004), .B0(n28751), .C0(n35855), .Y(
        n24005) );
  OAI211XL U28744 ( .A0(n30958), .A1(n24006), .B0(n24005), .C0(n34583), .Y(
        n15383) );
  INVXL U28745 ( .A(conv_1[154]), .Y(n24013) );
  AOI21XL U28746 ( .A0(n24009), .A1(n24008), .B0(n24007), .Y(n24011) );
  NAND2XL U28747 ( .A(conv_1[154]), .B(n24011), .Y(n24010) );
  OAI211XL U28748 ( .A0(conv_1[154]), .A1(n24011), .B0(n24499), .C0(n24010), 
        .Y(n24012) );
  OAI211XL U28749 ( .A0(n34048), .A1(n24013), .B0(n35489), .C0(n24012), .Y(
        n16309) );
  INVXL U28750 ( .A(conv_2[94]), .Y(n24020) );
  AOI21XL U28751 ( .A0(n24016), .A1(n24015), .B0(n24014), .Y(n24018) );
  NAND2XL U28752 ( .A(conv_2[94]), .B(n24018), .Y(n24017) );
  OAI211XL U28753 ( .A0(conv_2[94]), .A1(n24018), .B0(n32052), .C0(n24017), 
        .Y(n24019) );
  OAI211XL U28754 ( .A0(n34447), .A1(n24020), .B0(n34408), .C0(n24019), .Y(
        n15233) );
  ADDFXL U28755 ( .A(conv_3[242]), .B(n24023), .CI(n24022), .CO(n29658), .S(
        n23555) );
  AOI222XL U28756 ( .A0(n29657), .A1(n29658), .B0(n29657), .B1(conv_3[243]), 
        .C0(n29658), .C1(conv_3[243]), .Y(n24024) );
  INVXL U28757 ( .A(n24024), .Y(n24025) );
  NAND2XL U28758 ( .A(conv_3[244]), .B(n24028), .Y(n24027) );
  OAI211XL U28759 ( .A0(conv_3[244]), .A1(n24028), .B0(n35336), .C0(n24027), 
        .Y(n24029) );
  OAI211XL U28760 ( .A0(n35706), .A1(n24030), .B0(n34097), .C0(n24029), .Y(
        n15763) );
  AOI22XL U28761 ( .A0(n25299), .A1(conv_2[360]), .B0(n16673), .B1(conv_2[405]), .Y(n24032) );
  NAND2XL U28762 ( .A(n24032), .B(n24031), .Y(n24949) );
  INVXL U28763 ( .A(n24949), .Y(n25459) );
  AOI22XL U28764 ( .A0(n16666), .A1(conv_2[315]), .B0(n16662), .B1(conv_2[330]), .Y(n24034) );
  AOI22XL U28765 ( .A0(n25299), .A1(conv_2[300]), .B0(n16673), .B1(conv_2[345]), .Y(n24033) );
  NAND2XL U28766 ( .A(n24034), .B(n24033), .Y(n24948) );
  INVXL U28767 ( .A(n24948), .Y(n25464) );
  AOI222XL U28768 ( .A0(n34902), .A1(n36246), .B0(n22690), .B1(conv_2[420]), 
        .C0(n25306), .C1(conv_2[435]), .Y(n25458) );
  AOI22XL U28769 ( .A0(n16662), .A1(conv_2[150]), .B0(n16673), .B1(conv_2[165]), .Y(n24036) );
  AOI22XL U28770 ( .A0(n22762), .A1(conv_2[135]), .B0(n22690), .B1(conv_2[120]), .Y(n24035) );
  NAND2XL U28771 ( .A(n24036), .B(n24035), .Y(n34929) );
  INVXL U28772 ( .A(n34929), .Y(n24954) );
  OAI22XL U28773 ( .A0(n25458), .A1(n26474), .B0(n24954), .B1(n28479), .Y(
        n24051) );
  AOI22XL U28774 ( .A0(n16662), .A1(conv_2[210]), .B0(n16673), .B1(conv_2[225]), .Y(n24038) );
  AOI22XL U28775 ( .A0(n22762), .A1(conv_2[195]), .B0(n22690), .B1(conv_2[180]), .Y(n24037) );
  NAND2XL U28776 ( .A(n24038), .B(n24037), .Y(n25098) );
  INVXL U28777 ( .A(n25098), .Y(n34935) );
  INVXL U28778 ( .A(conv_2[285]), .Y(n34456) );
  AOI22XL U28779 ( .A0(n34984), .A1(n34932), .B0(n34931), .B1(n26451), .Y(
        n24049) );
  AOI22XL U28780 ( .A0(n16662), .A1(conv_2[90]), .B0(n18240), .B1(conv_2[105]), 
        .Y(n24045) );
  AOI22XL U28781 ( .A0(n22762), .A1(conv_2[75]), .B0(n18658), .B1(conv_2[60]), 
        .Y(n24044) );
  NAND2XL U28782 ( .A(n24045), .B(n24044), .Y(n34930) );
  AOI22XL U28783 ( .A0(n22762), .A1(conv_2[15]), .B0(n16673), .B1(conv_2[45]), 
        .Y(n24047) );
  AOI22XL U28784 ( .A0(n16662), .A1(conv_2[30]), .B0(n22690), .B1(conv_2[0]), 
        .Y(n24046) );
  NAND2XL U28785 ( .A(n24047), .B(n24046), .Y(n25100) );
  OAI211XL U28786 ( .A0(n34935), .A1(n28577), .B0(n24049), .C0(n24048), .Y(
        n24050) );
  AOI22XL U28787 ( .A0(n16670), .A1(n25199), .B0(n34984), .B1(n24778), .Y(
        n24055) );
  OAI22XL U28788 ( .A0(n25623), .A1(n28575), .B0(n34983), .B1(n25624), .Y(
        n24053) );
  OAI22XL U28789 ( .A0(n25620), .A1(n26474), .B0(n25030), .B1(n28479), .Y(
        n24052) );
  AOI211XL U28790 ( .A0(n28556), .A1(n25628), .B0(n24053), .C0(n24052), .Y(
        n24054) );
  OAI211XL U28791 ( .A0(n34989), .A1(n24783), .B0(n24055), .C0(n24054), .Y(
        n24133) );
  AOI22XL U28792 ( .A0(n28556), .A1(n25132), .B0(n25501), .B1(n24056), .Y(
        n24060) );
  OAI22XL U28793 ( .A0(n25502), .A1(n26473), .B0(n24982), .B1(n28479), .Y(
        n24058) );
  OAI22XL U28794 ( .A0(n24727), .A1(n35135), .B0(n34989), .B1(n24726), .Y(
        n24057) );
  NAND2XL U28795 ( .A(n24060), .B(n24059), .Y(n34878) );
  AOI22XL U28796 ( .A0(n16665), .A1(n24061), .B0(n25174), .B1(n26451), .Y(
        n24065) );
  INVXL U28797 ( .A(n25175), .Y(n25572) );
  OAI22XL U28798 ( .A0(n25574), .A1(n26473), .B0(n25572), .B1(n28479), .Y(
        n24063) );
  OAI22XL U28799 ( .A0(n25573), .A1(n26474), .B0(n25583), .B1(n28575), .Y(
        n24062) );
  AOI211XL U28800 ( .A0(n28556), .A1(n25571), .B0(n24063), .C0(n24062), .Y(
        n24064) );
  OAI211XL U28801 ( .A0(n34989), .A1(n24766), .B0(n24065), .C0(n24064), .Y(
        n24118) );
  INVXL U28802 ( .A(n25155), .Y(n25608) );
  AOI22XL U28803 ( .A0(n28528), .A1(n25600), .B0(n34984), .B1(n25608), .Y(
        n24069) );
  OAI22XL U28804 ( .A0(n25604), .A1(n28553), .B0(n25602), .B1(n34983), .Y(
        n24067) );
  OAI22XL U28805 ( .A0(n25154), .A1(n26474), .B0(n25603), .B1(n28577), .Y(
        n24066) );
  OAI211XL U28806 ( .A0(n34989), .A1(n24761), .B0(n24069), .C0(n24068), .Y(
        n24117) );
  INVXL U28807 ( .A(n25589), .Y(n24747) );
  OAI22XL U28808 ( .A0(n25586), .A1(n34983), .B0(n25590), .B1(n28553), .Y(
        n24071) );
  OAI22XL U28809 ( .A0(n25597), .A1(n28479), .B0(n25587), .B1(n28577), .Y(
        n24070) );
  AOI211XL U28810 ( .A0(n16671), .A1(n25183), .B0(n24071), .C0(n24070), .Y(
        n24072) );
  OAI211XL U28811 ( .A0(n34989), .A1(n24753), .B0(n24073), .C0(n24072), .Y(
        n24126) );
  NOR4XL U28812 ( .A(n34878), .B(n24118), .C(n24117), .D(n24126), .Y(n24092)
         );
  AOI22XL U28813 ( .A0(n34984), .A1(n24730), .B0(n25519), .B1(n26451), .Y(
        n24077) );
  OAI22XL U28814 ( .A0(n25141), .A1(n28577), .B0(n25513), .B1(n28479), .Y(
        n24075) );
  OAI22XL U28815 ( .A0(n25140), .A1(n26474), .B0(n25514), .B1(n28575), .Y(
        n24074) );
  AOI211XL U28816 ( .A0(n26470), .A1(n24735), .B0(n24075), .C0(n24074), .Y(
        n24076) );
  OAI211XL U28817 ( .A0(n25518), .A1(n28553), .B0(n24077), .C0(n24076), .Y(
        n24108) );
  INVXL U28818 ( .A(n25528), .Y(n24080) );
  INVXL U28819 ( .A(n25147), .Y(n25529) );
  OAI22XL U28820 ( .A0(n25527), .A1(n26473), .B0(n25529), .B1(n34983), .Y(
        n24079) );
  OAI22XL U28821 ( .A0(n25536), .A1(n26474), .B0(n25148), .B1(n28577), .Y(
        n24078) );
  AOI211XL U28822 ( .A0(n16659), .A1(n24080), .B0(n24079), .C0(n24078), .Y(
        n24081) );
  OAI211XL U28823 ( .A0(n34989), .A1(n24738), .B0(n24082), .C0(n24081), .Y(
        n24107) );
  INVXL U28824 ( .A(n25543), .Y(n24746) );
  AOI22XL U28825 ( .A0(n28556), .A1(n24746), .B0(n25542), .B1(n26451), .Y(
        n24086) );
  OAI22XL U28826 ( .A0(n25163), .A1(n26473), .B0(n25540), .B1(n28553), .Y(
        n24084) );
  OAI22XL U28827 ( .A0(n25550), .A1(n28575), .B0(n25541), .B1(n26474), .Y(
        n24083) );
  AOI211XL U28828 ( .A0(n28528), .A1(n25547), .B0(n24084), .C0(n24083), .Y(
        n24085) );
  OAI211XL U28829 ( .A0(n34989), .A1(n24743), .B0(n24086), .C0(n24085), .Y(
        n24106) );
  AOI22XL U28830 ( .A0(n28528), .A1(n25563), .B0(n25560), .B1(n26451), .Y(
        n24090) );
  OAI22XL U28831 ( .A0(n25566), .A1(n28577), .B0(n25556), .B1(n28575), .Y(
        n24088) );
  OAI22XL U28832 ( .A0(n25557), .A1(n26474), .B0(n25559), .B1(n26473), .Y(
        n24087) );
  AOI211XL U28833 ( .A0(n16665), .A1(n25558), .B0(n24088), .C0(n24087), .Y(
        n24089) );
  OAI211XL U28834 ( .A0(n34989), .A1(n24772), .B0(n24090), .C0(n24089), .Y(
        n24119) );
  NOR4XL U28835 ( .A(n24108), .B(n24107), .C(n24106), .D(n24119), .Y(n24091)
         );
  AOI21XL U28836 ( .A0(n24092), .A1(n24091), .B0(pool[59]), .Y(n24111) );
  OAI21XL U28837 ( .A0(n24962), .A1(n26409), .B0(n24093), .Y(n24095) );
  AOI222XL U28838 ( .A0(n25470), .A1(n36245), .B0(n25105), .B1(n22370), .C0(
        n24956), .C1(n28407), .Y(n24702) );
  OAI22XL U28839 ( .A0(n24702), .A1(n26575), .B0(n34989), .B1(n24704), .Y(
        n24094) );
  AOI211XL U28840 ( .A0(n28465), .A1(n24707), .B0(n24095), .C0(n24094), .Y(
        n24686) );
  AOI22XL U28841 ( .A0(n16667), .A1(n24715), .B0(n16670), .B1(n25127), .Y(
        n24099) );
  OAI22XL U28842 ( .A0(n25490), .A1(n26474), .B0(n25491), .B1(n26473), .Y(
        n24097) );
  OAI22XL U28843 ( .A0(n25119), .A1(n34983), .B0(n25124), .B1(n28575), .Y(
        n24096) );
  AOI211XL U28844 ( .A0(n34992), .A1(n25122), .B0(n24097), .C0(n24096), .Y(
        n24098) );
  OAI211XL U28845 ( .A0(n34989), .A1(n24716), .B0(n24099), .C0(n24098), .Y(
        n34876) );
  OAI22XL U28846 ( .A0(n24971), .A1(n19767), .B0(n25113), .B1(n28575), .Y(
        n24103) );
  AOI22XL U28847 ( .A0(n16667), .A1(n25115), .B0(n34984), .B1(n25487), .Y(
        n24101) );
  NAND2XL U28848 ( .A(n28465), .B(n24714), .Y(n24100) );
  OAI211XL U28849 ( .A0(n24708), .A1(n34989), .B0(n24101), .C0(n24100), .Y(
        n24102) );
  AOI211XL U28850 ( .A0(n28528), .A1(n25114), .B0(n24103), .C0(n24102), .Y(
        n34875) );
  AOI222XL U28851 ( .A0(n24136), .A1(pool[56]), .B0(n24136), .B1(n34875), .C0(
        pool[56]), .C1(n34875), .Y(n24104) );
  AOI222XL U28852 ( .A0(n34877), .A1(n34876), .B0(n34877), .B1(n24104), .C0(
        n34876), .C1(n24104), .Y(n24105) );
  AOI222XL U28853 ( .A0(pool[58]), .A1(n24686), .B0(pool[58]), .B1(n24105), 
        .C0(n24686), .C1(n24105), .Y(n24110) );
  NAND4XL U28854 ( .A(n34878), .B(n24108), .C(n24107), .D(n24106), .Y(n24109)
         );
  OAI22XL U28855 ( .A0(n25652), .A1(n34983), .B0(n25211), .B1(n26473), .Y(
        n24115) );
  AOI2BB2XL U28856 ( .B0(n16670), .B1(n25651), .A0N(n28577), .A1N(n25654), .Y(
        n24112) );
  OAI211XL U28857 ( .A0(n34989), .A1(n24793), .B0(n24113), .C0(n24112), .Y(
        n24114) );
  AOI211XL U28858 ( .A0(n16671), .A1(n25647), .B0(n24115), .C0(n24114), .Y(
        n24116) );
  INVXL U28859 ( .A(n24116), .Y(n24128) );
  AOI22XL U28860 ( .A0(n16667), .A1(n25632), .B0(n16670), .B1(n25643), .Y(
        n24124) );
  OAI22XL U28861 ( .A0(n25637), .A1(n26473), .B0(n25205), .B1(n28575), .Y(
        n24121) );
  OAI22XL U28862 ( .A0(n25636), .A1(n34983), .B0(n25634), .B1(n26474), .Y(
        n24120) );
  AOI211XL U28863 ( .A0(n26470), .A1(n24122), .B0(n24121), .C0(n24120), .Y(
        n24123) );
  OAI211XL U28864 ( .A0(n24125), .A1(n28479), .B0(n24124), .C0(n24123), .Y(
        n24129) );
  NAND4XL U28865 ( .A(pool[59]), .B(n24127), .C(n24126), .D(n24129), .Y(n24131) );
  NOR3XL U28866 ( .A(pool[59]), .B(n24129), .C(n24128), .Y(n24130) );
  NAND2XL U28867 ( .A(n34880), .B(pool[55]), .Y(n24135) );
  OAI21XL U28868 ( .A0(n24136), .A1(n34880), .B0(n24135), .Y(N29271) );
  INVXL U28869 ( .A(conv_1[180]), .Y(n24140) );
  OAI211XL U28870 ( .A0(n24138), .A1(conv_1[180]), .B0(n33778), .C0(n24137), 
        .Y(n24139) );
  OAI211XL U28871 ( .A0(n35368), .A1(n24140), .B0(n34773), .C0(n24139), .Y(
        n16283) );
  INVXL U28872 ( .A(conv_1[197]), .Y(n24146) );
  XOR2XL U28873 ( .A(n24142), .B(n24141), .Y(n24144) );
  NAND2XL U28874 ( .A(conv_1[197]), .B(n24144), .Y(n24143) );
  OAI211XL U28875 ( .A0(conv_1[197]), .A1(n24144), .B0(n24499), .C0(n24143), 
        .Y(n24145) );
  OAI211XL U28876 ( .A0(n35384), .A1(n24146), .B0(n33542), .C0(n24145), .Y(
        n16266) );
  INVXL U28877 ( .A(conv_1[181]), .Y(n24150) );
  OAI211XL U28878 ( .A0(n24148), .A1(conv_1[181]), .B0(n33778), .C0(n24147), 
        .Y(n24149) );
  OAI211XL U28879 ( .A0(n35368), .A1(n24150), .B0(n33067), .C0(n24149), .Y(
        n16282) );
  INVXL U28880 ( .A(conv_1[306]), .Y(n24157) );
  AOI21XL U28881 ( .A0(n24153), .A1(n28644), .B0(n24152), .Y(n24155) );
  NAND2XL U28882 ( .A(conv_1[306]), .B(n24155), .Y(n24154) );
  OAI211XL U28883 ( .A0(conv_1[306]), .A1(n24155), .B0(n30090), .C0(n24154), 
        .Y(n24156) );
  OAI211XL U28884 ( .A0(n33863), .A1(n24157), .B0(n34682), .C0(n24156), .Y(
        n16157) );
  INVXL U28885 ( .A(conv_1[313]), .Y(n24808) );
  NAND3XL U28886 ( .A(conv_1[312]), .B(n24175), .C(n24159), .Y(n24810) );
  OR3XL U28887 ( .A(n24175), .B(conv_1[312]), .C(n24159), .Y(n24809) );
  NAND2XL U28888 ( .A(n24810), .B(n24809), .Y(n24161) );
  NAND2XL U28889 ( .A(conv_1[313]), .B(n24161), .Y(n24160) );
  OAI211XL U28890 ( .A0(conv_1[313]), .A1(n24161), .B0(n34028), .C0(n24160), 
        .Y(n24162) );
  OAI211XL U28891 ( .A0(n33863), .A1(n24808), .B0(n16652), .C0(n24162), .Y(
        n16150) );
  OAI2BB1XL U28892 ( .A0N(n28644), .A1N(n28649), .B0(n24163), .Y(n24165) );
  NAND2XL U28893 ( .A(n24167), .B(n24165), .Y(n24164) );
  OAI211XL U28894 ( .A0(n24167), .A1(n24165), .B0(n24378), .C0(n24164), .Y(
        n24166) );
  OAI211XL U28895 ( .A0(n33863), .A1(n24167), .B0(n34544), .C0(n24166), .Y(
        n16154) );
  INVXL U28896 ( .A(conv_1[199]), .Y(n24173) );
  NAND2XL U28897 ( .A(conv_1[199]), .B(n24171), .Y(n24170) );
  OAI211XL U28898 ( .A0(conv_1[199]), .A1(n24171), .B0(n32611), .C0(n24170), 
        .Y(n24172) );
  OAI211XL U28899 ( .A0(n35384), .A1(n24173), .B0(n35489), .C0(n24172), .Y(
        n16264) );
  INVXL U28900 ( .A(conv_1[312]), .Y(n24179) );
  AOI21XL U28901 ( .A0(n24175), .A1(n28644), .B0(n24174), .Y(n24177) );
  NAND2XL U28902 ( .A(conv_1[312]), .B(n24177), .Y(n24176) );
  OAI211XL U28903 ( .A0(conv_1[312]), .A1(n24177), .B0(n33778), .C0(n24176), 
        .Y(n24178) );
  OAI211XL U28904 ( .A0(n33863), .A1(n24179), .B0(n34281), .C0(n24178), .Y(
        n16151) );
  INVXL U28905 ( .A(conv_2[300]), .Y(n24183) );
  OAI211XL U28906 ( .A0(n24181), .A1(conv_2[300]), .B0(n30090), .C0(n24180), 
        .Y(n24182) );
  OAI211XL U28907 ( .A0(n35976), .A1(n24183), .B0(n24182), .C0(n34583), .Y(
        n15363) );
  INVXL U28908 ( .A(conv_2[303]), .Y(n24189) );
  XOR2XL U28909 ( .A(n24185), .B(n24184), .Y(n24187) );
  NAND2XL U28910 ( .A(conv_2[303]), .B(n24187), .Y(n24186) );
  OAI211XL U28911 ( .A0(conv_2[303]), .A1(n24187), .B0(n34028), .C0(n24186), 
        .Y(n24188) );
  OAI211XL U28912 ( .A0(n35976), .A1(n24189), .B0(n24188), .C0(n34105), .Y(
        n15255) );
  INVXL U28913 ( .A(conv_2[349]), .Y(n24197) );
  AOI21XL U28914 ( .A0(n24193), .A1(n24192), .B0(n24191), .Y(n24195) );
  NAND2XL U28915 ( .A(conv_2[349]), .B(n24195), .Y(n24194) );
  OAI211XL U28916 ( .A0(conv_2[349]), .A1(n24195), .B0(n33788), .C0(n24194), 
        .Y(n24196) );
  OAI211XL U28917 ( .A0(n36010), .A1(n24197), .B0(n34408), .C0(n24196), .Y(
        n15216) );
  OAI211XL U28918 ( .A0(n24199), .A1(conv_2[15]), .B0(n32611), .C0(n24198), 
        .Y(n24200) );
  OAI211XL U28919 ( .A0(n30412), .A1(n24201), .B0(n34583), .C0(n24200), .Y(
        n15382) );
  INVXL U28920 ( .A(conv_3[378]), .Y(n24207) );
  NAND2XL U28921 ( .A(conv_3[378]), .B(n24205), .Y(n24204) );
  OAI211XL U28922 ( .A0(conv_3[378]), .A1(n24205), .B0(n32181), .C0(n24204), 
        .Y(n24206) );
  OAI211XL U28923 ( .A0(n34168), .A1(n24207), .B0(n35574), .C0(n24206), .Y(
        n15790) );
  INVXL U28924 ( .A(conv_2[419]), .Y(n33325) );
  NAND2XL U28925 ( .A(n24209), .B(conv_2[405]), .Y(n28069) );
  OAI211XL U28926 ( .A0(n24209), .A1(conv_2[405]), .B0(n32052), .C0(n28069), 
        .Y(n24210) );
  OAI211XL U28927 ( .A0(n36047), .A1(n24211), .B0(n24210), .C0(n34583), .Y(
        n15356) );
  INVXL U28928 ( .A(conv_2[16]), .Y(n24215) );
  OAI211XL U28929 ( .A0(n24213), .A1(conv_2[16]), .B0(n33982), .C0(n24212), 
        .Y(n24214) );
  OAI211XL U28930 ( .A0(n30412), .A1(n24215), .B0(n35847), .C0(n24214), .Y(
        n15346) );
  INVXL U28931 ( .A(conv_1[195]), .Y(n24219) );
  OAI211XL U28932 ( .A0(n24217), .A1(conv_1[195]), .B0(n33778), .C0(n24216), 
        .Y(n24218) );
  OAI211XL U28933 ( .A0(n35384), .A1(n24219), .B0(n34773), .C0(n24218), .Y(
        n16268) );
  INVXL U28934 ( .A(conv_1[196]), .Y(n24223) );
  OAI211XL U28935 ( .A0(n24221), .A1(conv_1[196]), .B0(n33778), .C0(n24220), 
        .Y(n24222) );
  OAI211XL U28936 ( .A0(n35384), .A1(n24223), .B0(n33067), .C0(n24222), .Y(
        n16267) );
  INVXL U28937 ( .A(conv_1[303]), .Y(n24229) );
  NAND2XL U28938 ( .A(conv_1[303]), .B(n24227), .Y(n24226) );
  OAI211XL U28939 ( .A0(conv_1[303]), .A1(n24227), .B0(n32052), .C0(n24226), 
        .Y(n24228) );
  OAI211XL U28940 ( .A0(n33863), .A1(n24229), .B0(n24228), .C0(n32867), .Y(
        n16160) );
  AOI22XL U28941 ( .A0(n24378), .A1(intadd_2_SUM_0_), .B0(conv_1[2]), .B1(
        n24536), .Y(n24230) );
  NAND2XL U28942 ( .A(n24230), .B(n33542), .Y(n16461) );
  AOI22XL U28943 ( .A0(n32656), .A1(n24234), .B0(conv_1[362]), .B1(n24233), 
        .Y(n24235) );
  NAND2XL U28944 ( .A(n24235), .B(n33542), .Y(n16101) );
  AOI22XL U28945 ( .A0(n32611), .A1(n24238), .B0(conv_3[62]), .B1(n32606), .Y(
        n24239) );
  NAND2XL U28946 ( .A(n24239), .B(n35566), .Y(n15847) );
  AOI22XL U28947 ( .A0(n32611), .A1(n24243), .B0(conv_1[334]), .B1(n24242), 
        .Y(n24244) );
  NAND2XL U28948 ( .A(n24244), .B(n35489), .Y(n16129) );
  AOI22XL U28949 ( .A0(n24378), .A1(intadd_2_SUM_2_), .B0(conv_1[4]), .B1(
        n24536), .Y(n24245) );
  NAND2XL U28950 ( .A(n24245), .B(n35489), .Y(n16459) );
  AOI22XL U28951 ( .A0(n32656), .A1(n24248), .B0(conv_3[377]), .B1(n32623), 
        .Y(n24249) );
  NAND2XL U28952 ( .A(n24249), .B(n35566), .Y(n15826) );
  ADDFX1 U28953 ( .A(conv_2[62]), .B(n24251), .CI(n24250), .CO(n26743), .S(
        n24252) );
  AOI22XL U28954 ( .A0(n32611), .A1(n24252), .B0(conv_2[62]), .B1(n33730), .Y(
        n24253) );
  NAND2XL U28955 ( .A(n24253), .B(n34621), .Y(n15307) );
  AOI22XL U28956 ( .A0(n32611), .A1(intadd_0_SUM_0_), .B0(conv_2[2]), .B1(
        n33566), .Y(n24254) );
  NAND2XL U28957 ( .A(n24254), .B(n34621), .Y(n15311) );
  AOI22XL U28958 ( .A0(n32656), .A1(n24257), .B0(conv_2[152]), .B1(n24358), 
        .Y(n24258) );
  NAND2XL U28959 ( .A(n24258), .B(n34621), .Y(n15301) );
  AOI21XL U28960 ( .A0(n24261), .A1(n24260), .B0(n24259), .Y(n24263) );
  NAND2XL U28961 ( .A(conv_3[454]), .B(n24263), .Y(n24262) );
  OAI211XL U28962 ( .A0(conv_3[454]), .A1(n24263), .B0(n36020), .C0(n24262), 
        .Y(n24264) );
  OAI211XL U28963 ( .A0(n35805), .A1(n24265), .B0(n34097), .C0(n24264), .Y(
        n15749) );
  OAI2BB1XL U28964 ( .A0N(n24270), .A1N(n24268), .B0(n24267), .Y(n24269) );
  OAI211XL U28965 ( .A0(n35865), .A1(n24270), .B0(n35847), .C0(n24269), .Y(
        n15345) );
  ADDFX1 U28966 ( .A(conv_1[243]), .B(n24272), .CI(n24271), .CO(n24440), .S(
        n24273) );
  AOI22XL U28967 ( .A0(n34028), .A1(n24273), .B0(conv_1[243]), .B1(n33658), 
        .Y(n24274) );
  NAND2XL U28968 ( .A(n24274), .B(n32867), .Y(n16220) );
  NAND2XL U28969 ( .A(n30672), .B(conv_1[345]), .Y(n24276) );
  OR2XL U28970 ( .A(n24276), .B(n26717), .Y(n34764) );
  INVXL U28971 ( .A(conv_1[346]), .Y(n24524) );
  NAND2XL U28972 ( .A(n35272), .B(n24276), .Y(n24275) );
  OAI211XL U28973 ( .A0(n35272), .A1(n24276), .B0(n34762), .C0(n24275), .Y(
        n24522) );
  OAI21XL U28974 ( .A0(n33403), .A1(n26717), .B0(n29761), .Y(n24278) );
  INVXL U28975 ( .A(n24278), .Y(n29762) );
  INVXL U28976 ( .A(conv_1[347]), .Y(n29767) );
  OAI22XL U28977 ( .A0(n33403), .A1(n29761), .B0(n29762), .B1(n29767), .Y(
        n24315) );
  AOI22XL U28978 ( .A0(n16657), .A1(n24280), .B0(conv_1[348]), .B1(n34763), 
        .Y(n24281) );
  NAND2XL U28979 ( .A(n24281), .B(n32867), .Y(n16115) );
  AOI22XL U28980 ( .A0(n28751), .A1(n24284), .B0(conv_1[153]), .B1(n24429), 
        .Y(n24285) );
  NAND2XL U28981 ( .A(n24285), .B(n32867), .Y(n16310) );
  AOI22XL U28982 ( .A0(n33822), .A1(n24289), .B0(conv_1[288]), .B1(n24288), 
        .Y(n24290) );
  NAND2XL U28983 ( .A(n24290), .B(n32867), .Y(n16175) );
  AOI22XL U28984 ( .A0(n33788), .A1(n24294), .B0(conv_1[213]), .B1(n24293), 
        .Y(n24295) );
  NAND2XL U28985 ( .A(n24295), .B(n32867), .Y(n16250) );
  ADDFX1 U28986 ( .A(conv_2[318]), .B(n24297), .CI(n24296), .CO(n23104), .S(
        n24299) );
  AOI22XL U28987 ( .A0(n36020), .A1(n24299), .B0(conv_2[318]), .B1(n24298), 
        .Y(n24300) );
  NAND2XL U28988 ( .A(n24300), .B(n34105), .Y(n15254) );
  AOI22XL U28989 ( .A0(n33778), .A1(n24304), .B0(conv_2[333]), .B1(n24303), 
        .Y(n24305) );
  NAND2XL U28990 ( .A(n24305), .B(n34105), .Y(n15253) );
  NAND2XL U28991 ( .A(conv_2[525]), .B(n28124), .Y(n24306) );
  OAI2BB1XL U28992 ( .A0N(n18913), .A1N(n24306), .B0(n34498), .Y(n29775) );
  NAND2XL U28993 ( .A(n34497), .B(n28126), .Y(n29776) );
  OAI21XL U28994 ( .A0(n29780), .A1(n29775), .B0(n29776), .Y(n24308) );
  NAND2XL U28995 ( .A(n35853), .B(n24308), .Y(n24307) );
  OAI31XL U28996 ( .A0(n35853), .A1(n33429), .A2(n24308), .B0(n24307), .Y(
        n27055) );
  NAND2XL U28997 ( .A(n24308), .B(n28128), .Y(n24309) );
  OAI2BB1XL U28998 ( .A0N(conv_2[527]), .A1N(n27055), .B0(n24309), .Y(n27684)
         );
  AOI22XL U28999 ( .A0(n32052), .A1(n24310), .B0(conv_2[528]), .B1(n33624), 
        .Y(n24311) );
  NAND2XL U29000 ( .A(n24311), .B(n34105), .Y(n15240) );
  AOI22XL U29001 ( .A0(n24378), .A1(n24313), .B0(conv_1[157]), .B1(n24429), 
        .Y(n24314) );
  NAND2XL U29002 ( .A(n24314), .B(n34682), .Y(n16306) );
  NOR2X1 U29003 ( .A(conv_1[351]), .B(n33643), .Y(n33644) );
  NOR2X1 U29004 ( .A(n33644), .B(n28847), .Y(n28809) );
  INVXL U29005 ( .A(conv_1[350]), .Y(n26367) );
  NOR2X1 U29006 ( .A(n26364), .B(n26367), .Y(n33645) );
  AOI21XL U29007 ( .A0(n33645), .A1(conv_1[351]), .B0(n35441), .Y(n28810) );
  AOI22XL U29008 ( .A0(n32660), .A1(n24320), .B0(conv_1[353]), .B1(n34763), 
        .Y(n24321) );
  NAND2XL U29009 ( .A(n24321), .B(n34696), .Y(n16110) );
  AOI22XL U29010 ( .A0(n34666), .A1(n24324), .B0(conv_3[213]), .B1(n35662), 
        .Y(n24325) );
  NAND2XL U29011 ( .A(n24325), .B(n35574), .Y(n15801) );
  ADDFX1 U29012 ( .A(conv_3[408]), .B(n24327), .CI(n24326), .CO(n26815), .S(
        n24328) );
  AOI22XL U29013 ( .A0(n27932), .A1(n24328), .B0(conv_3[408]), .B1(n32546), 
        .Y(n24329) );
  NAND2XL U29014 ( .A(n24329), .B(n35574), .Y(n15788) );
  ADDFX1 U29015 ( .A(conv_3[3]), .B(n24331), .CI(n24330), .CO(n24368), .S(
        n24332) );
  AOI22XL U29016 ( .A0(n36020), .A1(n24332), .B0(conv_3[3]), .B1(n27508), .Y(
        n24333) );
  NAND2XL U29017 ( .A(n24333), .B(n35574), .Y(n15815) );
  NAND2XL U29018 ( .A(conv_3[345]), .B(n27043), .Y(n27042) );
  OAI21XL U29019 ( .A0(n30536), .A1(n26717), .B0(n27042), .Y(n30569) );
  OAI21XL U29020 ( .A0(conv_3[346]), .A1(n30568), .B0(n30569), .Y(n30511) );
  OAI2BB1XL U29021 ( .A0N(n27619), .A1N(n34762), .B0(n30511), .Y(n24334) );
  INVXL U29022 ( .A(n24334), .Y(n30512) );
  INVXL U29023 ( .A(conv_3[347]), .Y(n30517) );
  OAI22XL U29024 ( .A0(n18997), .A1(n30511), .B0(n30512), .B1(n30517), .Y(
        n26715) );
  AOI22XL U29025 ( .A0(n28751), .A1(n24335), .B0(conv_3[348]), .B1(n33747), 
        .Y(n24336) );
  NAND2XL U29026 ( .A(n24336), .B(n35574), .Y(n15792) );
  AOI22XL U29027 ( .A0(n24499), .A1(n24339), .B0(conv_2[454]), .B1(n33606), 
        .Y(n24340) );
  NAND2XL U29028 ( .A(n24340), .B(n34408), .Y(n15209) );
  AOI22XL U29029 ( .A0(n33788), .A1(intadd_0_SUM_2_), .B0(conv_2[4]), .B1(
        n33566), .Y(n24341) );
  NAND2XL U29030 ( .A(n24341), .B(n34408), .Y(n15239) );
  INVXL U29031 ( .A(conv_1[82]), .Y(n34058) );
  OAI31XL U29032 ( .A0(conv_1[80]), .A1(n24931), .A2(conv_1[81]), .B0(n34053), 
        .Y(n34051) );
  OAI2BB1XL U29033 ( .A0N(n34058), .A1N(n34051), .B0(n34053), .Y(n24919) );
  AOI21XL U29034 ( .A0(n34052), .A1(conv_1[82]), .B0(n34053), .Y(n24920) );
  AOI22XL U29035 ( .A0(n32611), .A1(n24343), .B0(conv_1[84]), .B1(n24342), .Y(
        n24344) );
  NAND2XL U29036 ( .A(n24344), .B(n34281), .Y(n16379) );
  NAND2XL U29037 ( .A(n27230), .B(n34717), .Y(n24348) );
  ADDFX1 U29038 ( .A(conv_1[107]), .B(n24346), .CI(n24345), .CO(n31371), .S(
        n22934) );
  AOI222XL U29039 ( .A0(n31370), .A1(n31371), .B0(n31370), .B1(conv_1[108]), 
        .C0(n31371), .C1(conv_1[108]), .Y(n24347) );
  NAND2XL U29040 ( .A(n24348), .B(n24347), .Y(n32881) );
  INVXL U29041 ( .A(conv_1[110]), .Y(n29297) );
  AOI22XL U29042 ( .A0(n33778), .A1(n24350), .B0(conv_1[112]), .B1(n25090), 
        .Y(n24351) );
  NAND2XL U29043 ( .A(n24351), .B(n34696), .Y(n16351) );
  NOR2X1 U29044 ( .A(conv_2[126]), .B(n33803), .Y(n33804) );
  NOR2X1 U29045 ( .A(n33804), .B(n30443), .Y(n30061) );
  AOI21XL U29046 ( .A0(n33805), .A1(conv_2[126]), .B0(n34344), .Y(n30062) );
  AOI22XL U29047 ( .A0(n32611), .A1(n24355), .B0(conv_2[128]), .B1(n33801), 
        .Y(n24356) );
  NAND2XL U29048 ( .A(n24356), .B(n35859), .Y(n15120) );
  ADDFXL U29049 ( .A(conv_2[155]), .B(n34626), .CI(n24357), .CO(n24530), .S(
        n24359) );
  AOI22XL U29050 ( .A0(n24378), .A1(n24359), .B0(conv_2[155]), .B1(n24358), 
        .Y(n24360) );
  NAND2XL U29051 ( .A(n24360), .B(n35859), .Y(n15103) );
  INVXL U29052 ( .A(conv_2[131]), .Y(n34355) );
  OAI31XL U29053 ( .A0(conv_2[130]), .A1(conv_2[129]), .A2(n34343), .B0(n34344), .Y(n34350) );
  NAND2XL U29054 ( .A(conv_2[129]), .B(n34343), .Y(n30071) );
  AOI22XL U29055 ( .A0(n32611), .A1(n24362), .B0(conv_2[132]), .B1(n33801), 
        .Y(n24363) );
  NAND2XL U29056 ( .A(n24363), .B(n35859), .Y(n15116) );
  AOI22XL U29057 ( .A0(n32611), .A1(n24366), .B0(conv_3[530]), .B1(n33714), 
        .Y(n24367) );
  NAND2XL U29058 ( .A(n24367), .B(n35588), .Y(n15393) );
  NOR2X1 U29059 ( .A(conv_3[5]), .B(n28687), .Y(n24371) );
  INVXL U29060 ( .A(n28687), .Y(n24370) );
  INVXL U29061 ( .A(conv_3[5]), .Y(n28689) );
  INVXL U29062 ( .A(n31194), .Y(n24372) );
  INVXL U29063 ( .A(conv_3[8]), .Y(n31196) );
  OAI21XL U29064 ( .A0(conv_3[8]), .A1(n31194), .B0(n34379), .Y(n24373) );
  AOI22XL U29065 ( .A0(n24378), .A1(n24374), .B0(conv_3[10]), .B1(n27508), .Y(
        n24375) );
  NAND2XL U29066 ( .A(n24375), .B(n35588), .Y(n15738) );
  AOI22XL U29067 ( .A0(n24378), .A1(n24377), .B0(conv_3[7]), .B1(n27508), .Y(
        n24379) );
  NAND2XL U29068 ( .A(n24379), .B(n35588), .Y(n15741) );
  INVXL U29069 ( .A(pixel[49]), .Y(n24402) );
  INVXL U29070 ( .A(pixel[48]), .Y(n24381) );
  AOI22XL U29071 ( .A0(n22896), .A1(n24402), .B0(n24381), .B1(n23672), .Y(
        N17542) );
  INVXL U29072 ( .A(pixel[45]), .Y(n24389) );
  INVXL U29073 ( .A(pixel[44]), .Y(n24406) );
  AOI22XL U29074 ( .A0(n22896), .A1(n24389), .B0(n24406), .B1(n23672), .Y(
        N17538) );
  INVXL U29075 ( .A(pixel[51]), .Y(n24382) );
  INVXL U29076 ( .A(pixel[50]), .Y(n24403) );
  AOI22XL U29077 ( .A0(n22896), .A1(n24382), .B0(n24403), .B1(n23672), .Y(
        N17544) );
  INVXL U29078 ( .A(pixel[31]), .Y(n24399) );
  INVXL U29079 ( .A(pixel[30]), .Y(n24410) );
  AOI22XL U29080 ( .A0(n22896), .A1(n24399), .B0(n24410), .B1(n23672), .Y(
        N17524) );
  INVXL U29081 ( .A(pixel[38]), .Y(n24397) );
  INVXL U29082 ( .A(pixel[37]), .Y(n24392) );
  AOI22XL U29083 ( .A0(n22896), .A1(n24397), .B0(n24392), .B1(n23672), .Y(
        N17531) );
  INVXL U29084 ( .A(pixel[43]), .Y(n24405) );
  INVXL U29085 ( .A(pixel[42]), .Y(n24383) );
  AOI22XL U29086 ( .A0(n22896), .A1(n24405), .B0(n24383), .B1(n23672), .Y(
        N17536) );
  INVXL U29087 ( .A(pixel[47]), .Y(n24380) );
  INVXL U29088 ( .A(pixel[46]), .Y(n24390) );
  AOI22XL U29089 ( .A0(n22896), .A1(n24380), .B0(n24390), .B1(n23672), .Y(
        N17540) );
  AOI22XL U29090 ( .A0(n22896), .A1(n24381), .B0(n24380), .B1(n23672), .Y(
        N17541) );
  INVXL U29091 ( .A(pixel[36]), .Y(n24391) );
  INVXL U29092 ( .A(pixel[35]), .Y(n24388) );
  AOI22XL U29093 ( .A0(n22896), .A1(n24391), .B0(n24388), .B1(n23672), .Y(
        N17529) );
  INVXL U29094 ( .A(pixel[52]), .Y(n24508) );
  AOI22XL U29095 ( .A0(n22896), .A1(n24508), .B0(n24382), .B1(n23672), .Y(
        N17545) );
  INVXL U29096 ( .A(pixel[41]), .Y(n24395) );
  AOI22XL U29097 ( .A0(n22896), .A1(n24383), .B0(n24395), .B1(n23672), .Y(
        N17535) );
  NAND2XL U29098 ( .A(conv_1[242]), .B(n24385), .Y(n24384) );
  OAI211XL U29099 ( .A0(conv_1[242]), .A1(n24385), .B0(n32181), .C0(n24384), 
        .Y(n24386) );
  OAI211XL U29100 ( .A0(n35417), .A1(n24387), .B0(n24386), .C0(n33542), .Y(
        n16221) );
  INVXL U29101 ( .A(pixel[34]), .Y(n24393) );
  AOI22XL U29102 ( .A0(n22896), .A1(n24388), .B0(n24393), .B1(n23672), .Y(
        N17528) );
  AOI22XL U29103 ( .A0(n22896), .A1(n24390), .B0(n24389), .B1(n23672), .Y(
        N17539) );
  AOI22XL U29104 ( .A0(n22896), .A1(n24392), .B0(n24391), .B1(n23672), .Y(
        N17530) );
  INVXL U29105 ( .A(pixel[33]), .Y(n24394) );
  AOI22XL U29106 ( .A0(n22896), .A1(n24393), .B0(n24394), .B1(n23672), .Y(
        N17527) );
  INVXL U29107 ( .A(pixel[32]), .Y(n24400) );
  AOI22XL U29108 ( .A0(n22896), .A1(n24394), .B0(n24400), .B1(n23672), .Y(
        N17526) );
  INVXL U29109 ( .A(pixel[40]), .Y(n24396) );
  AOI22XL U29110 ( .A0(n22896), .A1(n24395), .B0(n24396), .B1(n23672), .Y(
        N17534) );
  INVXL U29111 ( .A(pixel[39]), .Y(n24398) );
  AOI22XL U29112 ( .A0(n22896), .A1(n24396), .B0(n24398), .B1(n23672), .Y(
        N17533) );
  AOI22XL U29113 ( .A0(n22896), .A1(n24398), .B0(n24397), .B1(n23672), .Y(
        N17532) );
  AOI22XL U29114 ( .A0(n22896), .A1(n24400), .B0(n24399), .B1(n23672), .Y(
        N17525) );
  INVXL U29115 ( .A(pixel[15]), .Y(n24404) );
  AOI22XL U29116 ( .A0(n22896), .A1(n24404), .B0(n24401), .B1(n23672), .Y(
        N17508) );
  AOI22XL U29117 ( .A0(n22896), .A1(n24403), .B0(n24402), .B1(n23672), .Y(
        N17543) );
  INVXL U29118 ( .A(pixel[16]), .Y(n24407) );
  AOI22XL U29119 ( .A0(n22896), .A1(n24407), .B0(n24404), .B1(n23672), .Y(
        N17509) );
  AOI22XL U29120 ( .A0(n22896), .A1(n24406), .B0(n24405), .B1(n23672), .Y(
        N17537) );
  INVXL U29121 ( .A(pixel[25]), .Y(n24420) );
  INVXL U29122 ( .A(pixel[24]), .Y(n24412) );
  AOI22XL U29123 ( .A0(n22896), .A1(n24420), .B0(n24412), .B1(n23672), .Y(
        N17518) );
  INVXL U29124 ( .A(pixel[19]), .Y(n24414) );
  INVXL U29125 ( .A(pixel[18]), .Y(n24409) );
  AOI22XL U29126 ( .A0(n22896), .A1(n24414), .B0(n24409), .B1(n23672), .Y(
        N17512) );
  INVXL U29127 ( .A(pixel[17]), .Y(n24408) );
  AOI22XL U29128 ( .A0(n22896), .A1(n24408), .B0(n24407), .B1(n23672), .Y(
        N17510) );
  AOI22XL U29129 ( .A0(n22896), .A1(n24409), .B0(n24408), .B1(n23672), .Y(
        N17511) );
  INVXL U29130 ( .A(pixel[29]), .Y(n24419) );
  AOI22XL U29131 ( .A0(n22896), .A1(n24410), .B0(n24419), .B1(n23672), .Y(
        N17523) );
  INVXL U29132 ( .A(pixel[23]), .Y(n24411) );
  INVXL U29133 ( .A(pixel[22]), .Y(n24417) );
  AOI22XL U29134 ( .A0(n22896), .A1(n24411), .B0(n24417), .B1(n23672), .Y(
        N17516) );
  AOI22XL U29135 ( .A0(n22896), .A1(n24412), .B0(n24411), .B1(n23672), .Y(
        N17517) );
  INVXL U29136 ( .A(pixel[27]), .Y(n24413) );
  INVXL U29137 ( .A(pixel[26]), .Y(n24421) );
  AOI22XL U29138 ( .A0(n22896), .A1(n24413), .B0(n24421), .B1(n23672), .Y(
        N17520) );
  INVXL U29139 ( .A(pixel[28]), .Y(n24418) );
  AOI22XL U29140 ( .A0(n22896), .A1(n24418), .B0(n24413), .B1(n23672), .Y(
        N17521) );
  INVXL U29141 ( .A(pixel[20]), .Y(n24415) );
  AOI22XL U29142 ( .A0(n22896), .A1(n24415), .B0(n24414), .B1(n23672), .Y(
        N17513) );
  INVXL U29143 ( .A(pixel[21]), .Y(n24416) );
  AOI22XL U29144 ( .A0(n22896), .A1(n24416), .B0(n24415), .B1(n23672), .Y(
        N17514) );
  AOI22XL U29145 ( .A0(n22896), .A1(n24417), .B0(n24416), .B1(n23672), .Y(
        N17515) );
  AOI22XL U29146 ( .A0(n22896), .A1(n24419), .B0(n24418), .B1(n23672), .Y(
        N17522) );
  AOI22XL U29147 ( .A0(n22896), .A1(n24421), .B0(n24420), .B1(n23672), .Y(
        N17519) );
  INVXL U29148 ( .A(filter_1[23]), .Y(n28218) );
  INVXL U29149 ( .A(filter_1[17]), .Y(n24423) );
  AOI22XL U29150 ( .A0(n36120), .A1(n28218), .B0(n24423), .B1(n28249), .Y(
        n14666) );
  INVXL U29151 ( .A(filter_1[53]), .Y(n24422) );
  AOI22XL U29152 ( .A0(n36120), .A1(n36151), .B0(n24422), .B1(n28249), .Y(
        n14672) );
  INVXL U29153 ( .A(filter_1[16]), .Y(n28216) );
  INVXL U29154 ( .A(filter_1[10]), .Y(n36119) );
  AOI22XL U29155 ( .A0(n36120), .A1(n28216), .B0(n36119), .B1(n28249), .Y(
        n14674) );
  INVXL U29156 ( .A(filter_1[47]), .Y(n24425) );
  AOI22XL U29157 ( .A0(n36120), .A1(n24422), .B0(n24425), .B1(n28249), .Y(
        n14671) );
  INVXL U29158 ( .A(filter_1[11]), .Y(n36121) );
  AOI22XL U29159 ( .A0(n36120), .A1(n24423), .B0(n36121), .B1(n28249), .Y(
        n14665) );
  INVXL U29160 ( .A(filter_1[48]), .Y(n28223) );
  AOI22XL U29161 ( .A0(n36120), .A1(n36124), .B0(n28223), .B1(n28249), .Y(
        n14717) );
  INVXL U29162 ( .A(filter_1[41]), .Y(n24424) );
  INVXL U29163 ( .A(filter_1[35]), .Y(n28227) );
  AOI22XL U29164 ( .A0(n36120), .A1(n24424), .B0(n28227), .B1(n28249), .Y(
        n14669) );
  AOI22XL U29165 ( .A0(n36120), .A1(n24425), .B0(n24424), .B1(n28249), .Y(
        n14670) );
  INVXL U29166 ( .A(filter_1[34]), .Y(n28231) );
  AOI22XL U29167 ( .A0(n36120), .A1(n24426), .B0(n28231), .B1(n28249), .Y(
        n14678) );
  ADDFX1 U29168 ( .A(conv_1[152]), .B(n24428), .CI(n24427), .CO(n24282), .S(
        n24430) );
  AOI22XL U29169 ( .A0(n33778), .A1(n24430), .B0(conv_1[152]), .B1(n24429), 
        .Y(n24431) );
  NAND2XL U29170 ( .A(n24431), .B(n33542), .Y(n16311) );
  NAND2XL U29171 ( .A(conv_1[241]), .B(n24435), .Y(n24434) );
  OAI211XL U29172 ( .A0(conv_1[241]), .A1(n24435), .B0(n33788), .C0(n24434), 
        .Y(n24436) );
  OAI211XL U29173 ( .A0(n35417), .A1(n24437), .B0(n24436), .C0(n33067), .Y(
        n16222) );
  INVXL U29174 ( .A(conv_1[244]), .Y(n24444) );
  AOI21XL U29175 ( .A0(n24440), .A1(n24439), .B0(n24438), .Y(n24442) );
  NAND2XL U29176 ( .A(conv_1[244]), .B(n24442), .Y(n24441) );
  OAI211XL U29177 ( .A0(conv_1[244]), .A1(n24442), .B0(n33778), .C0(n24441), 
        .Y(n24443) );
  OAI211XL U29178 ( .A0(n35417), .A1(n24444), .B0(n35489), .C0(n24443), .Y(
        n16219) );
  OAI21XL U29179 ( .A0(n18913), .A1(n32016), .B0(n24445), .Y(n30307) );
  AOI21XL U29180 ( .A0(conv_2[391]), .A1(n30307), .B0(n30306), .Y(n24447) );
  NAND2XL U29181 ( .A(n28128), .B(n27990), .Y(n24446) );
  AOI222XL U29182 ( .A0(n29056), .A1(n29055), .B0(n29056), .B1(conv_2[394]), 
        .C0(n29055), .C1(conv_2[394]), .Y(n24450) );
  NOR2X1 U29183 ( .A(n33953), .B(n24450), .Y(n28114) );
  AOI22XL U29184 ( .A0(n28751), .A1(n24452), .B0(conv_2[397]), .B1(n24451), 
        .Y(n24453) );
  NAND2XL U29185 ( .A(n24453), .B(n35859), .Y(n14941) );
  AOI22XL U29186 ( .A0(n33822), .A1(n24456), .B0(conv_2[367]), .B1(n24455), 
        .Y(n24457) );
  NAND2XL U29187 ( .A(n24457), .B(n35859), .Y(n14961) );
  AOI22XL U29188 ( .A0(n34028), .A1(n24460), .B0(conv_3[515]), .B1(n24479), 
        .Y(n24461) );
  NAND2XL U29189 ( .A(n24461), .B(n35588), .Y(n15403) );
  INVX1 U29190 ( .A(n33990), .Y(n33988) );
  NAND4XL U29191 ( .A(conv_3[30]), .B(n29680), .C(n29678), .D(n33990), .Y(
        n24463) );
  NAND2XL U29192 ( .A(conv_3[30]), .B(n29678), .Y(n24462) );
  INVXL U29193 ( .A(n24462), .Y(n33913) );
  AOI221XL U29194 ( .A0(n30536), .A1(n24462), .B0(n29680), .B1(n33913), .C0(
        n33988), .Y(n27528) );
  NAND2XL U29195 ( .A(n27528), .B(conv_3[31]), .Y(n27527) );
  NAND2XL U29196 ( .A(n24463), .B(n27527), .Y(n24464) );
  NAND2XL U29197 ( .A(n27619), .B(n24464), .Y(n30702) );
  AOI2BB1XL U29198 ( .A0N(n18997), .A1N(n33988), .B0(n24464), .Y(n24465) );
  INVXL U29199 ( .A(n24465), .Y(n30701) );
  NAND2XL U29200 ( .A(conv_3[32]), .B(n30701), .Y(n24466) );
  NAND2XL U29201 ( .A(n30702), .B(n24466), .Y(n29725) );
  AOI222XL U29202 ( .A0(n29726), .A1(conv_3[33]), .B0(n29726), .B1(n29725), 
        .C0(conv_3[33]), .C1(n29725), .Y(n24469) );
  NAND2XL U29203 ( .A(n24467), .B(n33990), .Y(n24468) );
  NAND2XL U29204 ( .A(n24469), .B(n24468), .Y(n29664) );
  NAND2XL U29205 ( .A(n35591), .B(n24470), .Y(n35584) );
  NAND2XL U29206 ( .A(conv_3[35]), .B(n35584), .Y(n31245) );
  NAND2XL U29207 ( .A(n33448), .B(conv_3[37]), .Y(n35590) );
  AOI21XL U29208 ( .A0(n31227), .A1(conv_3[39]), .B0(n33449), .Y(n31233) );
  INVXL U29209 ( .A(conv_3[44]), .Y(n31303) );
  AOI22XL U29210 ( .A0(n32611), .A1(n24471), .B0(conv_3[41]), .B1(n33444), .Y(
        n24472) );
  NAND2XL U29211 ( .A(n24472), .B(n35588), .Y(n15717) );
  NAND2XL U29212 ( .A(n31848), .B(n24475), .Y(n35647) );
  AOI21XL U29213 ( .A0(conv_3[200]), .A1(n35647), .B0(n35653), .Y(n31866) );
  AOI22XL U29214 ( .A0(n36020), .A1(n24476), .B0(conv_3[202]), .B1(n35655), 
        .Y(n24477) );
  NAND2XL U29215 ( .A(n24477), .B(n35588), .Y(n15611) );
  INVXL U29216 ( .A(conv_3[518]), .Y(n31184) );
  OAI31XL U29217 ( .A0(conv_3[516]), .A1(n31173), .A2(conv_3[517]), .B0(n31180), .Y(n31178) );
  INVXL U29218 ( .A(n31180), .Y(n31291) );
  AOI21XL U29219 ( .A0(n31184), .A1(n31178), .B0(n31291), .Y(n31147) );
  NAND2XL U29220 ( .A(conv_3[516]), .B(n31173), .Y(n31162) );
  AOI22XL U29221 ( .A0(n32656), .A1(n24480), .B0(conv_3[520]), .B1(n24479), 
        .Y(n24481) );
  NAND2XL U29222 ( .A(n24481), .B(n35588), .Y(n15398) );
  INVXL U29223 ( .A(conv_2[91]), .Y(n24485) );
  OAI211XL U29224 ( .A0(conv_2[91]), .A1(n24483), .B0(n33982), .C0(n24482), 
        .Y(n24484) );
  OAI211XL U29225 ( .A0(n34447), .A1(n24485), .B0(n24484), .C0(n35847), .Y(
        n15341) );
  OAI2BB1XL U29226 ( .A0N(n24488), .A1N(n24490), .B0(n24487), .Y(n24489) );
  OAI211XL U29227 ( .A0(n36010), .A1(n24490), .B0(n24489), .C0(n35847), .Y(
        n15324) );
  INVXL U29228 ( .A(conv_1[167]), .Y(n24494) );
  NAND2XL U29229 ( .A(conv_1[167]), .B(n24492), .Y(n24491) );
  OAI211XL U29230 ( .A0(conv_1[167]), .A1(n24492), .B0(n24499), .C0(n24491), 
        .Y(n24493) );
  OAI211XL U29231 ( .A0(n35346), .A1(n24494), .B0(n33542), .C0(n24493), .Y(
        n16296) );
  INVXL U29232 ( .A(conv_1[169]), .Y(n24502) );
  AOI21XL U29233 ( .A0(n24497), .A1(n24496), .B0(n24495), .Y(n24500) );
  NAND2XL U29234 ( .A(conv_1[169]), .B(n24500), .Y(n24498) );
  OAI211XL U29235 ( .A0(conv_1[169]), .A1(n24500), .B0(n24499), .C0(n24498), 
        .Y(n24501) );
  OAI211XL U29236 ( .A0(n35346), .A1(n24502), .B0(n35489), .C0(n24501), .Y(
        n16294) );
  INVXL U29237 ( .A(pixel[56]), .Y(n24506) );
  INVXL U29238 ( .A(pixel[55]), .Y(n24503) );
  AOI22XL U29239 ( .A0(n22896), .A1(n24506), .B0(n24503), .B1(n23672), .Y(
        N17549) );
  INVXL U29240 ( .A(pixel[54]), .Y(n24505) );
  AOI22XL U29241 ( .A0(n22896), .A1(n24503), .B0(n24505), .B1(n23672), .Y(
        N17548) );
  INVXL U29242 ( .A(pixel[59]), .Y(n24510) );
  INVXL U29243 ( .A(pixel[58]), .Y(n24504) );
  AOI22XL U29244 ( .A0(n22896), .A1(n24510), .B0(n24504), .B1(n23672), .Y(
        N17552) );
  INVXL U29245 ( .A(pixel[57]), .Y(n24507) );
  AOI22XL U29246 ( .A0(n22896), .A1(n24504), .B0(n24507), .B1(n23672), .Y(
        N17551) );
  INVXL U29247 ( .A(pixel[53]), .Y(n24509) );
  AOI22XL U29248 ( .A0(n22896), .A1(n24505), .B0(n24509), .B1(n23672), .Y(
        N17547) );
  AOI22XL U29249 ( .A0(n22896), .A1(n24507), .B0(n24506), .B1(n23672), .Y(
        N17550) );
  AOI22XL U29250 ( .A0(n22896), .A1(n24509), .B0(n24508), .B1(n23672), .Y(
        N17546) );
  INVXL U29251 ( .A(pixel[60]), .Y(n24511) );
  AOI22XL U29252 ( .A0(n22896), .A1(n24511), .B0(n24510), .B1(n23672), .Y(
        N17553) );
  INVXL U29253 ( .A(pixel[61]), .Y(n24512) );
  AOI22XL U29254 ( .A0(n22896), .A1(n24512), .B0(n24511), .B1(n23672), .Y(
        N17554) );
  INVXL U29255 ( .A(pixel[63]), .Y(n25087) );
  INVXL U29256 ( .A(pixel[62]), .Y(n24513) );
  AOI22XL U29257 ( .A0(n22896), .A1(n25087), .B0(n24513), .B1(n23672), .Y(
        N17556) );
  AOI22XL U29258 ( .A0(n22896), .A1(n24513), .B0(n24512), .B1(n23672), .Y(
        N17555) );
  INVXL U29259 ( .A(conv_1[302]), .Y(n24519) );
  NOR2BXL U29260 ( .AN(n24515), .B(n24514), .Y(n24517) );
  NAND2XL U29261 ( .A(conv_1[302]), .B(n24517), .Y(n24516) );
  OAI211XL U29262 ( .A0(conv_1[302]), .A1(n24517), .B0(n34028), .C0(n24516), 
        .Y(n24518) );
  OAI211XL U29263 ( .A0(n33863), .A1(n24519), .B0(n24518), .C0(n33542), .Y(
        n16161) );
  OAI2BB1XL U29264 ( .A0N(n24522), .A1N(n24524), .B0(n24521), .Y(n24523) );
  OAI211XL U29265 ( .A0(n35447), .A1(n24524), .B0(n24523), .C0(n33067), .Y(
        n16117) );
  OAI2BB1XL U29266 ( .A0N(n24529), .A1N(n24527), .B0(n24526), .Y(n24528) );
  OAI211XL U29267 ( .A0(n33863), .A1(n24529), .B0(n24528), .C0(n33067), .Y(
        n16162) );
  INVXL U29268 ( .A(n34626), .Y(n34623) );
  NAND2XL U29269 ( .A(conv_2[158]), .B(n29857), .Y(n28631) );
  NAND4XL U29270 ( .A(conv_2[161]), .B(conv_2[162]), .C(n34623), .D(n33946), 
        .Y(n26358) );
  INVXL U29271 ( .A(conv_2[162]), .Y(n33951) );
  INVXL U29272 ( .A(conv_2[161]), .Y(n33944) );
  NAND2XL U29273 ( .A(n34627), .B(n34625), .Y(n28635) );
  OAI21XL U29274 ( .A0(conv_2[160]), .A1(n28635), .B0(n34626), .Y(n33940) );
  NAND2XL U29275 ( .A(n33944), .B(n33940), .Y(n24531) );
  NAND3XL U29276 ( .A(n34626), .B(n33951), .C(n33947), .Y(n26357) );
  INVXL U29277 ( .A(conv_2[163]), .Y(n26361) );
  AOI22XL U29278 ( .A0(conv_2[163]), .A1(n26358), .B0(n26357), .B1(n26361), 
        .Y(n24533) );
  NAND2XL U29279 ( .A(conv_2[164]), .B(n24533), .Y(n24532) );
  OAI211XL U29280 ( .A0(conv_2[164]), .A1(n24533), .B0(n16657), .C0(n24532), 
        .Y(n24534) );
  OAI211XL U29281 ( .A0(n33853), .A1(n24535), .B0(n35859), .C0(n24534), .Y(
        n15094) );
  INVXL U29282 ( .A(conv_1[12]), .Y(n24542) );
  INVXL U29283 ( .A(n27278), .Y(n34547) );
  NOR2X1 U29284 ( .A(n27279), .B(conv_1[10]), .Y(n34548) );
  INVXL U29285 ( .A(n34548), .Y(n26298) );
  AOI32XL U29286 ( .A0(conv_1[11]), .A1(n34546), .A2(n34547), .B0(n24538), 
        .B1(n34546), .Y(n24540) );
  OAI2BB1XL U29287 ( .A0N(n24540), .A1N(n24542), .B0(n24539), .Y(n24541) );
  OAI211XL U29288 ( .A0(n34552), .A1(n24542), .B0(n34689), .C0(n24541), .Y(
        n16451) );
  MXI2XL U29289 ( .A(n24544), .B(n24543), .S0(n24570), .Y(n28209) );
  OAI2BB2XL U29290 ( .B0(n28210), .B1(n24546), .A0N(n24545), .A1N(n28209), .Y(
        n28208) );
  INVXL U29291 ( .A(affine_2[45]), .Y(n28207) );
  AOI22XL U29292 ( .A0(affine_2[45]), .A1(n33367), .B0(n16674), .B1(n24548), 
        .Y(n24549) );
  NAND2XL U29293 ( .A(n24549), .B(n33340), .Y(n16548) );
  OAI2BB1XL U29294 ( .A0N(n24552), .A1N(n24554), .B0(n24551), .Y(n24553) );
  OAI211XL U29295 ( .A0(n30994), .A1(n24554), .B0(n24553), .C0(n35847), .Y(
        n15329) );
  OAI2BB1XL U29296 ( .A0N(n24557), .A1N(n24559), .B0(n24556), .Y(n24558) );
  OAI211XL U29297 ( .A0(n35902), .A1(n24559), .B0(n24558), .C0(n35847), .Y(
        n15338) );
  MXI2XL U29298 ( .A(n24561), .B(n24560), .S0(n24570), .Y(n28396) );
  OAI2BB2XL U29299 ( .B0(n28397), .B1(n24563), .A0N(n24562), .A1N(n28396), .Y(
        n28395) );
  INVXL U29300 ( .A(affine_2[29]), .Y(n28394) );
  ADDFX1 U29301 ( .A(DP_OP_5170J1_126_4278_n26), .B(DP_OP_5170J1_126_4278_n28), 
        .CI(n24564), .CO(n28399), .S(n22090) );
  AOI22XL U29302 ( .A0(affine_2[29]), .A1(n33367), .B0(n16674), .B1(n24565), 
        .Y(n24566) );
  NAND2XL U29303 ( .A(n24566), .B(n33350), .Y(n16532) );
  AOI22XL U29304 ( .A0(n24569), .A1(n24568), .B0(n24567), .B1(n35018), .Y(
        N29333) );
  MXI2XL U29305 ( .A(n24571), .B(n18128), .S0(n24570), .Y(n28609) );
  OAI2BB2XL U29306 ( .B0(n28610), .B1(n24573), .A0N(n24572), .A1N(n28609), .Y(
        n28608) );
  INVXL U29307 ( .A(affine_2[13]), .Y(n28607) );
  ADDFX1 U29308 ( .A(DP_OP_5171J1_127_4278_n26), .B(DP_OP_5171J1_127_4278_n28), 
        .CI(n24574), .CO(n28612), .S(n22093) );
  AOI22XL U29309 ( .A0(affine_2[13]), .A1(n33367), .B0(n16674), .B1(n24575), 
        .Y(n24576) );
  NAND2XL U29310 ( .A(n24576), .B(n33368), .Y(n16566) );
  AOI22XL U29311 ( .A0(n36245), .A1(n28474), .B0(n24577), .B1(n28292), .Y(
        n26582) );
  INVXL U29312 ( .A(n26582), .Y(n24582) );
  OAI22XL U29313 ( .A0(n28470), .A1(n35184), .B0(n28469), .B1(n35200), .Y(
        n24581) );
  AOI2BB2XL U29314 ( .B0(n35236), .B1(n28475), .A0N(n35198), .A1N(n28472), .Y(
        n24579) );
  AOI22XL U29315 ( .A0(n35181), .A1(n28476), .B0(n35195), .B1(n28473), .Y(
        n24578) );
  OAI211XL U29316 ( .A0(n28471), .A1(n35196), .B0(n24579), .C0(n24578), .Y(
        n24580) );
  AOI211XL U29317 ( .A0(n28465), .A1(n24582), .B0(n24581), .C0(n24580), .Y(
        n24653) );
  OAI22XL U29318 ( .A0(n28518), .A1(n35196), .B0(n28516), .B1(n35200), .Y(
        n24586) );
  AOI22XL U29319 ( .A0(n36245), .A1(n28513), .B0(n28522), .B1(n28292), .Y(
        n26615) );
  INVXL U29320 ( .A(n28517), .Y(n26609) );
  AOI22XL U29321 ( .A0(n35195), .A1(n28512), .B0(n26609), .B1(n35207), .Y(
        n24584) );
  AOI2BB2XL U29322 ( .B0(n35236), .B1(n28514), .A0N(n35198), .A1N(n28519), .Y(
        n24583) );
  OAI211XL U29323 ( .A0(n35135), .A1(n26615), .B0(n24584), .C0(n24583), .Y(
        n24585) );
  AOI211XL U29324 ( .A0(n35181), .A1(n28515), .B0(n24586), .C0(n24585), .Y(
        n24652) );
  INVXL U29325 ( .A(n26569), .Y(n24589) );
  AOI22XL U29326 ( .A0(n35234), .A1(n26413), .B0(n26411), .B1(n35231), .Y(
        n24588) );
  AOI22XL U29327 ( .A0(n35236), .A1(n26570), .B0(n16660), .B1(n26412), .Y(
        n24587) );
  OAI211XL U29328 ( .A0(n24589), .A1(n35239), .B0(n24588), .C0(n24587), .Y(
        n24591) );
  AOI222XL U29329 ( .A0(n25335), .A1(n26374), .B0(n26411), .B1(n22369), .C0(
        n25334), .C1(n22362), .Y(n26573) );
  AOI22XL U29330 ( .A0(n36245), .A1(n25339), .B0(n25338), .B1(n28292), .Y(
        n26574) );
  OAI22XL U29331 ( .A0(n26573), .A1(n35159), .B0(n35135), .B1(n26574), .Y(
        n24590) );
  OAI22XL U29332 ( .A0(n28532), .A1(n35196), .B0(n28533), .B1(n35198), .Y(
        n24595) );
  AOI22XL U29333 ( .A0(n36245), .A1(n28537), .B0(n28527), .B1(n26374), .Y(
        n26626) );
  AOI2BB2XL U29334 ( .B0(n26444), .B1(n35207), .A0N(n35200), .A1N(n28531), .Y(
        n24593) );
  AOI22XL U29335 ( .A0(n35181), .A1(n28526), .B0(n35195), .B1(n28529), .Y(
        n24592) );
  OAI211XL U29336 ( .A0(n35135), .A1(n26626), .B0(n24593), .C0(n24592), .Y(
        n24594) );
  AOI211XL U29337 ( .A0(n35236), .A1(n28530), .B0(n24595), .C0(n24594), .Y(
        n24651) );
  NAND4XL U29338 ( .A(n24653), .B(n24652), .C(n24666), .D(n24651), .Y(n24634)
         );
  INVXL U29339 ( .A(pool[44]), .Y(n24667) );
  AOI22XL U29340 ( .A0(n36245), .A1(n28442), .B0(n28443), .B1(n26374), .Y(
        n26606) );
  OAI22XL U29341 ( .A0(n28439), .A1(n35196), .B0(n28440), .B1(n18208), .Y(
        n24599) );
  AOI22XL U29342 ( .A0(n16660), .A1(n28437), .B0(n16664), .B1(n25345), .Y(
        n24597) );
  AOI2BB2XL U29343 ( .B0(n28436), .B1(n35207), .A0N(n35239), .A1N(n28438), .Y(
        n24596) );
  OAI211XL U29344 ( .A0(n28449), .A1(n35202), .B0(n24597), .C0(n24596), .Y(
        n24598) );
  AOI211XL U29345 ( .A0(n28465), .A1(n26606), .B0(n24599), .C0(n24598), .Y(
        n24658) );
  OAI22XL U29346 ( .A0(n28503), .A1(n35202), .B0(n28511), .B1(n35184), .Y(
        n24603) );
  AOI22XL U29347 ( .A0(n35236), .A1(n28498), .B0(n35234), .B1(n26588), .Y(
        n24601) );
  INVXL U29348 ( .A(n28502), .Y(n26587) );
  INVXL U29349 ( .A(n28501), .Y(n26423) );
  AOI22XL U29350 ( .A0(n16660), .A1(n26587), .B0(n16664), .B1(n26423), .Y(
        n24600) );
  OAI211XL U29351 ( .A0(n28505), .A1(n35239), .B0(n24601), .C0(n24600), .Y(
        n24602) );
  AOI211XL U29352 ( .A0(n28465), .A1(n26593), .B0(n24603), .C0(n24602), .Y(
        n24657) );
  AOI22XL U29353 ( .A0(n36245), .A1(n28454), .B0(n28452), .B1(n28292), .Y(
        n26618) );
  OAI22XL U29354 ( .A0(n28457), .A1(n35239), .B0(n28456), .B1(n35198), .Y(
        n24608) );
  AOI22XL U29355 ( .A0(n35236), .A1(n28451), .B0(n35234), .B1(n26449), .Y(
        n24606) );
  AOI22XL U29356 ( .A0(n16664), .A1(n24604), .B0(n28450), .B1(n35207), .Y(
        n24605) );
  OAI211XL U29357 ( .A0(n28463), .A1(n35202), .B0(n24606), .C0(n24605), .Y(
        n24607) );
  AOI211XL U29358 ( .A0(n28465), .A1(n26618), .B0(n24608), .C0(n24607), .Y(
        n24650) );
  AOI22XL U29359 ( .A0(n36245), .A1(n28484), .B0(n28485), .B1(n26374), .Y(
        n26598) );
  INVXL U29360 ( .A(n26598), .Y(n26421) );
  OAI22XL U29361 ( .A0(n28489), .A1(n35198), .B0(n28491), .B1(n35202), .Y(
        n24612) );
  AOI22XL U29362 ( .A0(n35195), .A1(n28486), .B0(n35234), .B1(n26594), .Y(
        n24610) );
  AOI22XL U29363 ( .A0(n35236), .A1(n28487), .B0(n28494), .B1(n35207), .Y(
        n24609) );
  OAI211XL U29364 ( .A0(n28488), .A1(n35200), .B0(n24610), .C0(n24609), .Y(
        n24611) );
  AOI211XL U29365 ( .A0(n28465), .A1(n26421), .B0(n24612), .C0(n24611), .Y(
        n24654) );
  NAND4XL U29366 ( .A(n24658), .B(n24657), .C(n24650), .D(n24654), .Y(n24633)
         );
  AOI22XL U29367 ( .A0(n35195), .A1(n26537), .B0(n35236), .B1(n26538), .Y(
        n24614) );
  AOI22XL U29368 ( .A0(n16660), .A1(n26385), .B0(n26384), .B1(n35231), .Y(
        n24613) );
  OAI211XL U29369 ( .A0(n25376), .A1(n35196), .B0(n24614), .C0(n24613), .Y(
        n24617) );
  AOI222XL U29370 ( .A0(n24615), .A1(n26374), .B0(n26384), .B1(n22369), .C0(
        n25374), .C1(n22362), .Y(n26541) );
  AOI22XL U29371 ( .A0(n36245), .A1(n25378), .B0(n25380), .B1(n28292), .Y(
        n26542) );
  OAI22XL U29372 ( .A0(n26541), .A1(n35159), .B0(n35135), .B1(n26542), .Y(
        n24616) );
  INVXL U29373 ( .A(pool[42]), .Y(n34859) );
  OAI22XL U29374 ( .A0(n24618), .A1(n35143), .B0(n26555), .B1(n35198), .Y(
        n24621) );
  INVXL U29375 ( .A(n26401), .Y(n24619) );
  AOI222XL U29376 ( .A0(n26398), .A1(n28291), .B0(n24619), .B1(n28290), .C0(
        n26562), .C1(n28289), .Y(n26558) );
  OAI22XL U29377 ( .A0(N18471), .A1(n26558), .B0(n26557), .B1(n35135), .Y(
        n24620) );
  AOI211XL U29378 ( .A0(n35236), .A1(n26563), .B0(n24621), .C0(n24620), .Y(
        n24623) );
  NAND2XL U29379 ( .A(n35195), .B(n26399), .Y(n24622) );
  OAI211XL U29380 ( .A0(n26566), .A1(n35196), .B0(n24623), .C0(n24622), .Y(
        n34858) );
  INVXL U29381 ( .A(n25394), .Y(n24625) );
  AOI222XL U29382 ( .A0(n24625), .A1(n28292), .B0(n25400), .B1(n22369), .C0(
        n25392), .C1(n22362), .Y(n26550) );
  AOI22XL U29383 ( .A0(n35195), .A1(n26546), .B0(n35236), .B1(n26547), .Y(
        n24627) );
  AOI22XL U29384 ( .A0(n16660), .A1(n26395), .B0(n25400), .B1(n35231), .Y(
        n24626) );
  OAI211XL U29385 ( .A0(n26393), .A1(n35196), .B0(n24627), .C0(n24626), .Y(
        n24628) );
  AOI211XL U29386 ( .A0(n26554), .A1(n28465), .B0(n24629), .C0(n24628), .Y(
        n34857) );
  AOI222XL U29387 ( .A0(pool[40]), .A1(pool[41]), .B0(pool[40]), .B1(n34857), 
        .C0(pool[41]), .C1(n34857), .Y(n24630) );
  AOI222XL U29388 ( .A0(n34859), .A1(n34858), .B0(n34859), .B1(n24630), .C0(
        n34858), .C1(n24630), .Y(n24631) );
  AOI222XL U29389 ( .A0(n34862), .A1(pool[43]), .B0(n34862), .B1(n24631), .C0(
        pool[43]), .C1(n24631), .Y(n24632) );
  AOI221XL U29390 ( .A0(n24634), .A1(n24667), .B0(n24633), .B1(n24667), .C0(
        n24632), .Y(n24664) );
  AOI22XL U29391 ( .A0(n35181), .A1(n28410), .B0(n18197), .B1(n26632), .Y(
        n24638) );
  OAI2BB2XL U29392 ( .B0(n28415), .B1(n35200), .A0N(n28412), .A1N(n35195), .Y(
        n24636) );
  INVXL U29393 ( .A(n28413), .Y(n26462) );
  OAI22XL U29394 ( .A0(n35184), .A1(n26633), .B0(n26462), .B1(n35196), .Y(
        n24635) );
  AOI211XL U29395 ( .A0(n35236), .A1(n25312), .B0(n24636), .C0(n24635), .Y(
        n24637) );
  AOI22XL U29396 ( .A0(n36245), .A1(n28555), .B0(n28557), .B1(n26374), .Y(
        n26652) );
  AOI22XL U29397 ( .A0(n35195), .A1(n28558), .B0(n35236), .B1(n28560), .Y(
        n24643) );
  OAI22XL U29398 ( .A0(n28549), .A1(n35200), .B0(n28552), .B1(n35202), .Y(
        n24640) );
  OAI22XL U29399 ( .A0(n28563), .A1(n35196), .B0(n28550), .B1(n35184), .Y(
        n24639) );
  AOI211XL U29400 ( .A0(n16660), .A1(n24641), .B0(n24640), .C0(n24639), .Y(
        n24642) );
  OAI211XL U29401 ( .A0(n35135), .A1(n26652), .B0(n24643), .C0(n24642), .Y(
        n24659) );
  AOI22XL U29402 ( .A0(n36245), .A1(n24644), .B0(n28572), .B1(n28292), .Y(
        n26647) );
  AOI22XL U29403 ( .A0(n16660), .A1(n28583), .B0(n28570), .B1(n35207), .Y(
        n24648) );
  OAI22XL U29404 ( .A0(n26641), .A1(n35202), .B0(n28579), .B1(n35239), .Y(
        n24646) );
  OAI22XL U29405 ( .A0(n28580), .A1(n35200), .B0(n28576), .B1(n35196), .Y(
        n24645) );
  AOI211XL U29406 ( .A0(n35236), .A1(n28573), .B0(n24646), .C0(n24645), .Y(
        n24647) );
  OAI211XL U29407 ( .A0(n35135), .A1(n26647), .B0(n24648), .C0(n24647), .Y(
        n24649) );
  NOR3XL U29408 ( .A(pool[44]), .B(n24659), .C(n24649), .Y(n24662) );
  NAND2BXL U29409 ( .AN(n24650), .B(n24649), .Y(n24656) );
  OR4XL U29410 ( .A(n24654), .B(n24653), .C(n24652), .D(n24651), .Y(n24655) );
  NOR4XL U29411 ( .A(n24658), .B(n24657), .C(n24656), .D(n24655), .Y(n24660)
         );
  NAND4BXL U29412 ( .AN(n24666), .B(pool[44]), .C(n24660), .D(n24659), .Y(
        n24661) );
  AOI22XL U29413 ( .A0(n34860), .A1(n24667), .B0(n24666), .B1(n34861), .Y(
        N29260) );
  OAI2BB1XL U29414 ( .A0N(n24670), .A1N(n24672), .B0(n24669), .Y(n24671) );
  OAI211XL U29415 ( .A0(n35610), .A1(n24672), .B0(n24671), .C0(n33550), .Y(
        n15882) );
  INVXL U29416 ( .A(conv_1[44]), .Y(n33127) );
  NAND2XL U29417 ( .A(conv_1[30]), .B(n30672), .Y(n33433) );
  NAND2XL U29418 ( .A(n35272), .B(n33433), .Y(n24674) );
  OAI211XL U29419 ( .A0(n35272), .A1(n33433), .B0(n33990), .C0(n24674), .Y(
        n24676) );
  NOR2X1 U29420 ( .A(n24676), .B(n24678), .Y(n25073) );
  OAI2BB1XL U29421 ( .A0N(n24678), .A1N(n24676), .B0(n24675), .Y(n24677) );
  OAI211XL U29422 ( .A0(n35302), .A1(n24678), .B0(n24677), .C0(n33067), .Y(
        n16432) );
  NAND2XL U29423 ( .A(n24680), .B(n24679), .Y(n24682) );
  AOI211XL U29424 ( .A0(n24684), .A1(n24682), .B0(n36042), .C0(n24681), .Y(
        n24683) );
  AOI2BB1XL U29425 ( .A0N(n24684), .A1N(n35395), .B0(n24683), .Y(n24685) );
  NAND2XL U29426 ( .A(n24685), .B(n34544), .Y(n16245) );
  INVXL U29427 ( .A(n34880), .Y(n34874) );
  AOI22XL U29428 ( .A0(n34880), .A1(n24687), .B0(n24686), .B1(n34874), .Y(
        N29274) );
  NAND2XL U29429 ( .A(n27230), .B(n34422), .Y(n24692) );
  INVXL U29430 ( .A(n24688), .Y(n24689) );
  OAI21XL U29431 ( .A0(conv_1[258]), .A1(n24690), .B0(n24689), .Y(n24691) );
  OAI21XL U29432 ( .A0(n24695), .A1(n16655), .B0(n34080), .Y(n24694) );
  NAND2XL U29433 ( .A(n24696), .B(n34544), .Y(n16203) );
  INVXL U29434 ( .A(n25458), .Y(n24697) );
  AOI222XL U29435 ( .A0(n25100), .A1(n28291), .B0(n24697), .B1(n28290), .C0(
        n34931), .C1(n28289), .Y(n34928) );
  INVXL U29436 ( .A(n28304), .Y(n26561) );
  AOI22XL U29437 ( .A0(n16663), .A1(n34932), .B0(n34931), .B1(n26561), .Y(
        n24698) );
  OAI211XL U29438 ( .A0(n24954), .A1(n28553), .B0(n24699), .C0(n24698), .Y(
        n24700) );
  AOI22XL U29439 ( .A0(n16665), .A1(n25104), .B0(n28366), .B1(n25108), .Y(
        n24703) );
  OR2XL U29440 ( .A(n35241), .B(n25109), .Y(n25473) );
  OAI211XL U29441 ( .A0(n24704), .A1(n16701), .B0(n24703), .C0(n25473), .Y(
        n24705) );
  AOI22XL U29442 ( .A0(n28366), .A1(n24709), .B0(n16663), .B1(n25487), .Y(
        n24711) );
  OAI211XL U29443 ( .A0(n24971), .A1(n28304), .B0(n24711), .C0(n24710), .Y(
        n24712) );
  AOI222XL U29444 ( .A0(n24807), .A1(pool[61]), .B0(n24807), .B1(n34881), .C0(
        pool[61]), .C1(n34881), .Y(n24722) );
  AOI22XL U29445 ( .A0(n16665), .A1(n25122), .B0(n25496), .B1(n26561), .Y(
        n24721) );
  OAI22XL U29446 ( .A0(n25491), .A1(n28349), .B0(n25124), .B1(n26621), .Y(
        n24719) );
  OAI22XL U29447 ( .A0(n24717), .A1(n28467), .B0(n16701), .B1(n24716), .Y(
        n24718) );
  OAI211XL U29448 ( .A0(n25120), .A1(n28575), .B0(n24721), .C0(n24720), .Y(
        n34882) );
  INVXL U29449 ( .A(pool[62]), .Y(n34883) );
  AOI222XL U29450 ( .A0(n24722), .A1(n34882), .B0(n24722), .B1(n34883), .C0(
        n34882), .C1(n34883), .Y(n24723) );
  AOI222XL U29451 ( .A0(pool[63]), .A1(n34886), .B0(pool[63]), .B1(n24723), 
        .C0(n34886), .C1(n24723), .Y(n24777) );
  INVXL U29452 ( .A(pool[64]), .Y(n26151) );
  AOI22XL U29453 ( .A0(n16665), .A1(n25131), .B0(n25501), .B1(n26561), .Y(
        n24724) );
  OAI211XL U29454 ( .A0(n25502), .A1(n28349), .B0(n24725), .C0(n24724), .Y(
        n24729) );
  OAI22XL U29455 ( .A0(n24727), .A1(n34989), .B0(n16701), .B1(n24726), .Y(
        n24728) );
  OAI22XL U29456 ( .A0(n25518), .A1(n16672), .B0(n25514), .B1(n26621), .Y(
        n24734) );
  INVXL U29457 ( .A(n25141), .Y(n25517) );
  AOI22XL U29458 ( .A0(n34961), .A1(n25516), .B0(n16663), .B1(n24730), .Y(
        n24731) );
  OAI211XL U29459 ( .A0(n25513), .A1(n28553), .B0(n24732), .C0(n24731), .Y(
        n24733) );
  AOI211XL U29460 ( .A0(n34827), .A1(n24735), .B0(n24734), .C0(n24733), .Y(
        n24756) );
  OAI22XL U29461 ( .A0(n25527), .A1(n28349), .B0(n25528), .B1(n28553), .Y(
        n24740) );
  AOI2BB2XL U29462 ( .B0(n18463), .B1(n25531), .A0N(n18196), .A1N(n25536), .Y(
        n24737) );
  INVXL U29463 ( .A(n25148), .Y(n25530) );
  OAI211XL U29464 ( .A0(n26575), .A1(n24738), .B0(n24737), .C0(n24736), .Y(
        n24739) );
  AOI211XL U29465 ( .A0(n28324), .A1(n25526), .B0(n24740), .C0(n24739), .Y(
        n24755) );
  OAI22XL U29466 ( .A0(n25541), .A1(n18196), .B0(n25540), .B1(n16672), .Y(
        n24745) );
  AOI22XL U29467 ( .A0(n28366), .A1(n25162), .B0(n25542), .B1(n28372), .Y(
        n24742) );
  INVXL U29468 ( .A(n25163), .Y(n25544) );
  AOI22XL U29469 ( .A0(n16665), .A1(n25547), .B0(n16663), .B1(n25544), .Y(
        n24741) );
  OAI211XL U29470 ( .A0(n26575), .A1(n24743), .B0(n24742), .C0(n24741), .Y(
        n24744) );
  AOI22XL U29471 ( .A0(n16665), .A1(n24748), .B0(n16663), .B1(n24747), .Y(
        n24752) );
  INVXL U29472 ( .A(n25183), .Y(n25591) );
  OAI22XL U29473 ( .A0(n25591), .A1(n18196), .B0(n25587), .B1(n28575), .Y(
        n24750) );
  INVXL U29474 ( .A(n28372), .Y(n28333) );
  OAI22XL U29475 ( .A0(n25586), .A1(n28333), .B0(n25590), .B1(n16672), .Y(
        n24749) );
  AOI211XL U29476 ( .A0(n28324), .A1(n25588), .B0(n24750), .C0(n24749), .Y(
        n24751) );
  OAI211XL U29477 ( .A0(n26575), .A1(n24753), .B0(n24752), .C0(n24751), .Y(
        n24795) );
  NAND4BXL U29478 ( .AN(n24795), .B(n24756), .C(n24755), .D(n24754), .Y(n24774) );
  AOI22XL U29479 ( .A0(n34961), .A1(n25598), .B0(n25156), .B1(n28372), .Y(
        n24760) );
  OAI22XL U29480 ( .A0(n25603), .A1(n28575), .B0(n25604), .B1(n16672), .Y(
        n24758) );
  OAI2BB2XL U29481 ( .B0(n25155), .B1(n28349), .A0N(n25601), .A1N(n28324), .Y(
        n24757) );
  AOI211XL U29482 ( .A0(n16665), .A1(n25600), .B0(n24758), .C0(n24757), .Y(
        n24759) );
  OAI211XL U29483 ( .A0(n26575), .A1(n24761), .B0(n24760), .C0(n24759), .Y(
        n24799) );
  AOI2BB2XL U29484 ( .B0(n25174), .B1(n28372), .A0N(n26621), .A1N(n25583), .Y(
        n24765) );
  OAI22XL U29485 ( .A0(n25573), .A1(n18196), .B0(n25176), .B1(n34981), .Y(
        n24763) );
  OAI22XL U29486 ( .A0(n25575), .A1(n16672), .B0(n25574), .B1(n28349), .Y(
        n24762) );
  AOI211XL U29487 ( .A0(n16665), .A1(n25175), .B0(n24763), .C0(n24762), .Y(
        n24764) );
  OAI211XL U29488 ( .A0(n26575), .A1(n24766), .B0(n24765), .C0(n24764), .Y(
        n24798) );
  AOI22XL U29489 ( .A0(n34961), .A1(n25010), .B0(n28559), .B1(n25558), .Y(
        n24771) );
  OAI22XL U29490 ( .A0(n25566), .A1(n28575), .B0(n25556), .B1(n26621), .Y(
        n24769) );
  OAI22XL U29491 ( .A0(n25559), .A1(n28349), .B0(n24767), .B1(n28333), .Y(
        n24768) );
  AOI211XL U29492 ( .A0(n16670), .A1(n25563), .B0(n24769), .C0(n24768), .Y(
        n24770) );
  OAI211XL U29493 ( .A0(n26575), .A1(n24772), .B0(n24771), .C0(n24770), .Y(
        n24796) );
  NOR4BXL U29494 ( .AN(n26150), .B(n24799), .C(n24798), .D(n24796), .Y(n24773)
         );
  NAND2BXL U29495 ( .AN(n24774), .B(n24773), .Y(n24775) );
  AOI22XL U29496 ( .A0(n16665), .A1(n25619), .B0(n16663), .B1(n24778), .Y(
        n24782) );
  OAI22XL U29497 ( .A0(n25623), .A1(n26621), .B0(n28333), .B1(n25624), .Y(
        n24780) );
  INVXL U29498 ( .A(n25199), .Y(n25625) );
  OAI22XL U29499 ( .A0(n25620), .A1(n18196), .B0(n25625), .B1(n16672), .Y(
        n24779) );
  OAI22XL U29500 ( .A0(n25637), .A1(n28349), .B0(n25205), .B1(n26621), .Y(
        n24785) );
  OAI22XL U29501 ( .A0(n25634), .A1(n18196), .B0(n25636), .B1(n28333), .Y(
        n24784) );
  AOI211XL U29502 ( .A0(n18463), .A1(n25643), .B0(n24785), .C0(n24784), .Y(
        n24786) );
  OAI211XL U29503 ( .A0(n26575), .A1(n24788), .B0(n24787), .C0(n24786), .Y(
        n24794) );
  AOI22XL U29504 ( .A0(n34961), .A1(n25647), .B0(n16670), .B1(n25648), .Y(
        n24792) );
  OAI2BB2XL U29505 ( .B0(n25652), .B1(n28333), .A0N(n25657), .A1N(n28324), .Y(
        n24790) );
  OAI22XL U29506 ( .A0(n25211), .A1(n28349), .B0(n25654), .B1(n34981), .Y(
        n24789) );
  AOI211XL U29507 ( .A0(n18463), .A1(n25651), .B0(n24790), .C0(n24789), .Y(
        n24791) );
  OAI211XL U29508 ( .A0(n26575), .A1(n24793), .B0(n24792), .C0(n24791), .Y(
        n24797) );
  NOR3XL U29509 ( .A(pool[64]), .B(n24794), .C(n24797), .Y(n24802) );
  NAND4XL U29510 ( .A(n24800), .B(n24799), .C(n24798), .D(n24797), .Y(n24801)
         );
  NAND2XL U29511 ( .A(n34884), .B(pool[60]), .Y(n24806) );
  OAI21XL U29512 ( .A0(n24807), .A1(n34884), .B0(n24806), .Y(N29276) );
  AOI22XL U29513 ( .A0(conv_1[313]), .A1(n24810), .B0(n24809), .B1(n24808), 
        .Y(n24812) );
  NAND2XL U29514 ( .A(conv_1[314]), .B(n24812), .Y(n24811) );
  OAI211XL U29515 ( .A0(conv_1[314]), .A1(n24812), .B0(n32052), .C0(n24811), 
        .Y(n24813) );
  OAI211XL U29516 ( .A0(n33442), .A1(n24814), .B0(n34696), .C0(n24813), .Y(
        n16149) );
  OAI22XL U29517 ( .A0(n35178), .A1(n28553), .B0(n35170), .B1(n26473), .Y(
        n24818) );
  AOI22XL U29518 ( .A0(n16659), .A1(n28264), .B0(n28556), .B1(n35167), .Y(
        n24815) );
  OAI211XL U29519 ( .A0(n35171), .A1(n26474), .B0(n24816), .C0(n24815), .Y(
        n24817) );
  AOI22XL U29520 ( .A0(n36245), .A1(n26214), .B0(n26215), .B1(n26374), .Y(
        n35097) );
  INVXL U29521 ( .A(n28315), .Y(n35093) );
  AOI22XL U29522 ( .A0(n16665), .A1(n35094), .B0(n34984), .B1(n35093), .Y(
        n24822) );
  INVXL U29523 ( .A(n35100), .Y(n28316) );
  OAI22XL U29524 ( .A0(n34983), .A1(n35090), .B0(n28316), .B1(n28577), .Y(
        n24820) );
  OAI22XL U29525 ( .A0(n26213), .A1(n28575), .B0(n35089), .B1(n26474), .Y(
        n24819) );
  AOI211XL U29526 ( .A0(n34992), .A1(n35091), .B0(n24820), .C0(n24819), .Y(
        n24821) );
  OAI211XL U29527 ( .A0(n34989), .A1(n35097), .B0(n24822), .C0(n24821), .Y(
        n24893) );
  AOI22XL U29528 ( .A0(n36245), .A1(n26237), .B0(n26240), .B1(n28292), .Y(
        n35064) );
  INVXL U29529 ( .A(n35057), .Y(n28350) );
  INVXL U29530 ( .A(n28351), .Y(n35058) );
  OAI22XL U29531 ( .A0(n35056), .A1(n26474), .B0(n35058), .B1(n28479), .Y(
        n24824) );
  OAI22XL U29532 ( .A0(n35053), .A1(n26473), .B0(n35055), .B1(n28553), .Y(
        n24823) );
  AOI211XL U29533 ( .A0(n16667), .A1(n28350), .B0(n24824), .C0(n24823), .Y(
        n24825) );
  OAI211XL U29534 ( .A0(n34989), .A1(n35064), .B0(n24826), .C0(n24825), .Y(
        n24898) );
  INVXL U29535 ( .A(n24827), .Y(n35101) );
  OAI22XL U29536 ( .A0(n19767), .A1(n24828), .B0(n35103), .B1(n26473), .Y(
        n24831) );
  INVXL U29537 ( .A(n25770), .Y(n24829) );
  AOI222XL U29538 ( .A0(n24829), .A1(n28292), .B0(n35104), .B1(n22369), .C0(
        n26208), .C1(n22362), .Y(n35109) );
  OAI22XL U29539 ( .A0(n35109), .A1(n35135), .B0(n34989), .B1(n35108), .Y(
        n24830) );
  AOI211XL U29540 ( .A0(n16667), .A1(n35101), .B0(n24831), .C0(n24830), .Y(
        n24833) );
  NAND2XL U29541 ( .A(n28528), .B(n35102), .Y(n24832) );
  OAI211XL U29542 ( .A0(n35107), .A1(n28575), .B0(n24833), .C0(n24832), .Y(
        n24890) );
  AOI22XL U29543 ( .A0(n36245), .A1(n26191), .B0(n26192), .B1(n26374), .Y(
        n35049) );
  AOI22XL U29544 ( .A0(n28414), .A1(n35052), .B0(n26451), .B1(n35045), .Y(
        n24837) );
  INVXL U29545 ( .A(n25748), .Y(n35043) );
  OAI22XL U29546 ( .A0(n35042), .A1(n28553), .B0(n35041), .B1(n28479), .Y(
        n24835) );
  OAI22XL U29547 ( .A0(n28310), .A1(n28577), .B0(n26190), .B1(n26473), .Y(
        n24834) );
  AOI211XL U29548 ( .A0(n16671), .A1(n35043), .B0(n24835), .C0(n24834), .Y(
        n24836) );
  OAI211XL U29549 ( .A0(n34989), .A1(n35049), .B0(n24837), .C0(n24836), .Y(
        n24897) );
  INVXL U29550 ( .A(n26182), .Y(n35141) );
  OAI22XL U29551 ( .A0(n35141), .A1(n28577), .B0(n28276), .B1(n26473), .Y(
        n24841) );
  AOI22XL U29552 ( .A0(n36245), .A1(n25716), .B0(n25717), .B1(n28292), .Y(
        n35144) );
  AOI22XL U29553 ( .A0(n16659), .A1(n35140), .B0(n26451), .B1(n28278), .Y(
        n24839) );
  OAI211XL U29554 ( .A0(n34989), .A1(n35144), .B0(n24839), .C0(n24838), .Y(
        n24840) );
  AOI211XL U29555 ( .A0(n16665), .A1(n28280), .B0(n24841), .C0(n24840), .Y(
        n34998) );
  INVXL U29556 ( .A(pool[100]), .Y(n34993) );
  INVXL U29557 ( .A(n25712), .Y(n24842) );
  AOI222XL U29558 ( .A0(n24842), .A1(n26374), .B0(n35153), .B1(n22369), .C0(
        n26179), .C1(n22362), .Y(n35160) );
  AOI22XL U29559 ( .A0(n36245), .A1(n25715), .B0(n25707), .B1(n26374), .Y(
        n35158) );
  OAI22XL U29560 ( .A0(n35160), .A1(n35135), .B0(n34989), .B1(n35158), .Y(
        n24843) );
  AOI211XL U29561 ( .A0(n16667), .A1(n35151), .B0(n24844), .C0(n24843), .Y(
        n24845) );
  OAI211XL U29562 ( .A0(n19767), .A1(n28301), .B0(n24846), .C0(n24845), .Y(
        n34995) );
  AOI222XL U29563 ( .A0(n34993), .A1(n34996), .B0(n34993), .B1(n34995), .C0(
        n34996), .C1(n34995), .Y(n24847) );
  AOI222XL U29564 ( .A0(pool[102]), .A1(n34998), .B0(pool[102]), .B1(n24847), 
        .C0(n34998), .C1(n24847), .Y(n24854) );
  AOI22XL U29565 ( .A0(n28528), .A1(n35127), .B0(n34954), .B1(n26171), .Y(
        n24853) );
  INVXL U29566 ( .A(n25697), .Y(n24850) );
  AOI222XL U29567 ( .A0(n24850), .A1(n28292), .B0(n26171), .B1(n22369), .C0(
        n26170), .C1(n22362), .Y(n35136) );
  AOI22XL U29568 ( .A0(n36245), .A1(n25699), .B0(n25700), .B1(n28292), .Y(
        n35134) );
  OAI22XL U29569 ( .A0(n35136), .A1(n35135), .B0(n34989), .B1(n35134), .Y(
        n24851) );
  OAI211XL U29570 ( .A0(n35126), .A1(n28575), .B0(n24853), .C0(n24852), .Y(
        n34999) );
  INVXL U29571 ( .A(pool[103]), .Y(n35000) );
  AOI22XL U29572 ( .A0(n36245), .A1(n26200), .B0(n26199), .B1(n26374), .Y(
        n35076) );
  AOI2BB2X1 U29573 ( .B0(n34963), .B1(n35073), .A0N(n28479), .A1N(n35067), .Y(
        n24858) );
  OAI22XL U29574 ( .A0(n28321), .A1(n26474), .B0(n35065), .B1(n26473), .Y(
        n24856) );
  OAI22XL U29575 ( .A0(n34983), .A1(n35070), .B0(n35068), .B1(n28553), .Y(
        n24855) );
  AOI211XL U29576 ( .A0(n16667), .A1(n35069), .B0(n24856), .C0(n24855), .Y(
        n24857) );
  OAI211XL U29577 ( .A0(n26479), .A1(n35076), .B0(n24858), .C0(n24857), .Y(
        n24888) );
  AOI2BB2XL U29578 ( .B0(n26232), .B1(n28292), .A0N(n26374), .A1N(n26229), .Y(
        n35120) );
  AOI22XL U29579 ( .A0(n28414), .A1(n35115), .B0(n34984), .B1(n35116), .Y(
        n24863) );
  OAI22XL U29580 ( .A0(n34983), .A1(n24859), .B0(n35113), .B1(n28577), .Y(
        n24861) );
  OAI22XL U29581 ( .A0(n28339), .A1(n28479), .B0(n35112), .B1(n26474), .Y(
        n24860) );
  AOI211XL U29582 ( .A0(n16665), .A1(n35123), .B0(n24861), .C0(n24860), .Y(
        n24862) );
  OAI211XL U29583 ( .A0(n34989), .A1(n35120), .B0(n24863), .C0(n24862), .Y(
        n24887) );
  AOI22XL U29584 ( .A0(n16659), .A1(n35079), .B0(n16670), .B1(n35080), .Y(
        n24868) );
  AOI22XL U29585 ( .A0(n36245), .A1(n26223), .B0(n24864), .B1(n28292), .Y(
        n35088) );
  OAI22XL U29586 ( .A0(n35085), .A1(n28577), .B0(n35077), .B1(n26473), .Y(
        n24866) );
  OAI22XL U29587 ( .A0(n34983), .A1(n35081), .B0(n28332), .B1(n28575), .Y(
        n24865) );
  AOI211XL U29588 ( .A0(n26470), .A1(n35088), .B0(n24866), .C0(n24865), .Y(
        n24867) );
  OAI211XL U29589 ( .A0(n35078), .A1(n26474), .B0(n24868), .C0(n24867), .Y(
        n24886) );
  AOI22XL U29590 ( .A0(n36245), .A1(n26244), .B0(n26245), .B1(n26374), .Y(
        n35037) );
  AOI22XL U29591 ( .A0(n16659), .A1(n28344), .B0(n26451), .B1(n35034), .Y(
        n24872) );
  OAI22XL U29592 ( .A0(n35030), .A1(n26473), .B0(n26246), .B1(n28553), .Y(
        n24870) );
  OAI22XL U29593 ( .A0(n25732), .A1(n26474), .B0(n35033), .B1(n28577), .Y(
        n24869) );
  OAI211XL U29594 ( .A0(n34989), .A1(n35037), .B0(n24872), .C0(n24871), .Y(
        n24892) );
  NOR4XL U29595 ( .A(n24888), .B(n24887), .C(n24886), .D(n24892), .Y(n24873)
         );
  OAI22XL U29596 ( .A0(n35186), .A1(n26473), .B0(n35182), .B1(n26474), .Y(
        n24880) );
  AOI22XL U29597 ( .A0(n36245), .A1(n24876), .B0(n26275), .B1(n28292), .Y(
        n35192) );
  AOI22XL U29598 ( .A0(n28528), .A1(n35189), .B0(n26451), .B1(n28364), .Y(
        n24878) );
  OAI211XL U29599 ( .A0(n34989), .A1(n35192), .B0(n24878), .C0(n24877), .Y(
        n24879) );
  AOI211XL U29600 ( .A0(n16665), .A1(n35180), .B0(n24880), .C0(n24879), .Y(
        n24891) );
  OAI22XL U29601 ( .A0(n35201), .A1(n26474), .B0(n24881), .B1(n34981), .Y(
        n24885) );
  AOI22XL U29602 ( .A0(n36245), .A1(n26261), .B0(n26259), .B1(n26374), .Y(
        n35210) );
  AOI22XL U29603 ( .A0(n34984), .A1(n28373), .B0(n26451), .B1(n35206), .Y(
        n24883) );
  AOI22XL U29604 ( .A0(n16659), .A1(n35193), .B0(n16670), .B1(n28371), .Y(
        n24882) );
  OAI211XL U29605 ( .A0(n34989), .A1(n35210), .B0(n24883), .C0(n24882), .Y(
        n24884) );
  AOI211XL U29606 ( .A0(n16667), .A1(n28374), .B0(n24885), .C0(n24884), .Y(
        n24889) );
  INVXL U29607 ( .A(pool[104]), .Y(n24905) );
  NAND3XL U29608 ( .A(n24891), .B(n24889), .C(n24905), .Y(n24900) );
  NAND4BXL U29609 ( .AN(n24889), .B(n24888), .C(n24887), .D(n24886), .Y(n24896) );
  INVXL U29610 ( .A(n24890), .Y(n24904) );
  NAND4XL U29611 ( .A(pool[104]), .B(n24894), .C(n24893), .D(n24892), .Y(
        n24895) );
  INVXL U29612 ( .A(n35001), .Y(n34997) );
  AOI22XL U29613 ( .A0(n35001), .A1(n24905), .B0(n24904), .B1(n34997), .Y(
        N29320) );
  INVXL U29614 ( .A(conv_1[524]), .Y(n29250) );
  NAND4XL U29615 ( .A(conv_1[510]), .B(n27429), .C(n30672), .D(n34019), .Y(
        n24907) );
  NAND2XL U29616 ( .A(conv_1[510]), .B(n30672), .Y(n24906) );
  INVXL U29617 ( .A(n24906), .Y(n34017) );
  AOI221XL U29618 ( .A0(n35272), .A1(n24906), .B0(n27429), .B1(n34017), .C0(
        n27764), .Y(n27017) );
  NAND2XL U29619 ( .A(conv_1[511]), .B(n27017), .Y(n27016) );
  NAND2XL U29620 ( .A(n24907), .B(n27016), .Y(n24910) );
  NAND2XL U29621 ( .A(n33403), .B(n24910), .Y(n24908) );
  OAI31XL U29622 ( .A0(n33403), .A1(n27764), .A2(n24910), .B0(n24908), .Y(
        n26983) );
  NAND2XL U29623 ( .A(n24910), .B(n24909), .Y(n24911) );
  OAI2BB1XL U29624 ( .A0N(conv_1[512]), .A1N(n26983), .B0(n24911), .Y(n30455)
         );
  INVXL U29625 ( .A(n30267), .Y(n29246) );
  OAI21XL U29626 ( .A0(conv_1[516]), .A1(n27266), .B0(n29246), .Y(n25259) );
  NAND2XL U29627 ( .A(n25259), .B(n25258), .Y(n24915) );
  AOI211XL U29628 ( .A0(n24917), .A1(n24915), .B0(n36042), .C0(n24914), .Y(
        n24916) );
  AOI2BB1XL U29629 ( .A0N(n24917), .A1N(n35547), .B0(n24916), .Y(n24918) );
  NAND2XL U29630 ( .A(n24918), .B(n34682), .Y(n15946) );
  NAND2BXL U29631 ( .AN(n24920), .B(n24919), .Y(n24922) );
  AOI211XL U29632 ( .A0(n24924), .A1(n24922), .B0(n36042), .C0(n24921), .Y(
        n24923) );
  AOI2BB1XL U29633 ( .A0N(n24924), .A1N(n34057), .B0(n24923), .Y(n24925) );
  NAND2XL U29634 ( .A(n24925), .B(n34281), .Y(n16380) );
  OAI2BB1XL U29635 ( .A0N(conv_1[85]), .A1N(n26724), .B0(n26735), .Y(n26734)
         );
  AOI32XL U29636 ( .A0(conv_1[86]), .A1(n26735), .A2(n26734), .B0(n34053), 
        .B1(n26737), .Y(n24928) );
  AOI211XL U29637 ( .A0(n26736), .A1(n24928), .B0(n36042), .C0(n24927), .Y(
        n24929) );
  AOI2BB1XL U29638 ( .A0N(n26736), .A1N(n34057), .B0(n24929), .Y(n24930) );
  NAND2XL U29639 ( .A(n24930), .B(n34281), .Y(n16376) );
  AOI22XL U29640 ( .A0(n34053), .A1(n24932), .B0(n24931), .B1(n26735), .Y(
        n24934) );
  AOI211XL U29641 ( .A0(n24936), .A1(n24934), .B0(n36042), .C0(n24933), .Y(
        n24935) );
  AOI2BB1XL U29642 ( .A0N(n24936), .A1N(n34057), .B0(n24935), .Y(n24937) );
  NAND2XL U29643 ( .A(n24937), .B(n34281), .Y(n16383) );
  INVXL U29644 ( .A(conv_1[494]), .Y(n33358) );
  INVXL U29645 ( .A(conv_1[481]), .Y(n24942) );
  NAND2XL U29646 ( .A(n30672), .B(conv_1[480]), .Y(n27212) );
  NAND2XL U29647 ( .A(n35272), .B(n27212), .Y(n24938) );
  OAI211XL U29648 ( .A0(n35272), .A1(n27212), .B0(n33530), .C0(n24938), .Y(
        n24940) );
  OAI2BB1XL U29649 ( .A0N(n24942), .A1N(n24940), .B0(n24939), .Y(n24941) );
  OAI211XL U29650 ( .A0(n35544), .A1(n24942), .B0(n33067), .C0(n24941), .Y(
        n15982) );
  OAI2BB1XL U29651 ( .A0N(n24947), .A1N(n24945), .B0(n24944), .Y(n24946) );
  OAI211XL U29652 ( .A0(n33427), .A1(n24947), .B0(n33067), .C0(n24946), .Y(
        n15967) );
  AOI22XL U29653 ( .A0(n36244), .A1(n34931), .B0(n28289), .B1(n24948), .Y(
        n24951) );
  AOI22XL U29654 ( .A0(n25337), .A1(n34932), .B0(n25399), .B1(n24949), .Y(
        n24950) );
  OAI211XL U29655 ( .A0(n25458), .A1(n25393), .B0(n24951), .C0(n24950), .Y(
        n25103) );
  AOI22XL U29656 ( .A0(n26263), .A1(n25098), .B0(n26172), .B1(n34931), .Y(
        n24953) );
  OAI211XL U29657 ( .A0(n24954), .A1(n28577), .B0(n24953), .C0(n24952), .Y(
        n24955) );
  AOI22XL U29658 ( .A0(n25336), .A1(n25469), .B0(n25399), .B1(n25467), .Y(
        n24958) );
  AOI22XL U29659 ( .A0(n36244), .A1(n24956), .B0(n28289), .B1(n25468), .Y(
        n24957) );
  OAI211XL U29660 ( .A0(n24959), .A1(n25402), .B0(n24958), .C0(n24957), .Y(
        n25111) );
  AOI22XL U29661 ( .A0(n26263), .A1(n25105), .B0(n28528), .B1(n25108), .Y(
        n24960) );
  OAI211XL U29662 ( .A0(n24962), .A1(n26207), .B0(n24961), .C0(n24960), .Y(
        n24963) );
  OAI2BB2XL U29663 ( .B0(n25119), .B1(n16721), .A0N(n25489), .A1N(n28289), .Y(
        n24965) );
  OAI22XL U29664 ( .A0(n25491), .A1(n25402), .B0(n25490), .B1(n25393), .Y(
        n24964) );
  OAI22XL U29665 ( .A0(n25119), .A1(n26207), .B0(n25120), .B1(n16661), .Y(
        n24967) );
  OAI2BB2XL U29666 ( .B0(n25124), .B1(n28479), .A0N(n25122), .A1N(n16667), .Y(
        n24966) );
  OAI22XL U29667 ( .A0(n24971), .A1(n26207), .B0(n25113), .B1(n28479), .Y(
        n24975) );
  AOI2BB2XL U29668 ( .B0(n25337), .B1(n25487), .A0N(n25393), .A1N(n25477), .Y(
        n24970) );
  AOI22XL U29669 ( .A0(n25399), .A1(n25478), .B0(n28289), .B1(n25479), .Y(
        n24969) );
  OAI211XL U29670 ( .A0(n24971), .A1(n16721), .B0(n24970), .C0(n24969), .Y(
        n25118) );
  OAI2BB1XL U29671 ( .A0N(N18471), .A1N(n25118), .B0(n24973), .Y(n24974) );
  AOI222XL U29672 ( .A0(pool[46]), .A1(n34863), .B0(pool[46]), .B1(n25061), 
        .C0(n34863), .C1(n25061), .Y(n24976) );
  AOI222XL U29673 ( .A0(n34867), .A1(n34865), .B0(n34867), .B1(n24976), .C0(
        n34865), .C1(n24976), .Y(n24977) );
  AOI222XL U29674 ( .A0(pool[48]), .A1(n25446), .B0(pool[48]), .B1(n24977), 
        .C0(n25446), .C1(n24977), .Y(n25029) );
  AOI22XL U29675 ( .A0(n36244), .A1(n25501), .B0(n25399), .B1(n25503), .Y(
        n24979) );
  AOI22XL U29676 ( .A0(n25336), .A1(n25511), .B0(n28289), .B1(n25504), .Y(
        n24978) );
  OAI211XL U29677 ( .A0(n25502), .A1(n25402), .B0(n24979), .C0(n24978), .Y(
        n25138) );
  AOI22XL U29678 ( .A0(n26263), .A1(n25132), .B0(n28528), .B1(n25135), .Y(
        n24981) );
  OAI211XL U29679 ( .A0(n24982), .A1(n28577), .B0(n24981), .C0(n24980), .Y(
        n24983) );
  AOI21XL U29680 ( .A0(N18471), .A1(n25138), .B0(n24983), .Y(n25444) );
  OAI22XL U29681 ( .A0(n25527), .A1(n26285), .B0(n25536), .B1(n26274), .Y(
        n24988) );
  OAI22XL U29682 ( .A0(n25148), .A1(n16661), .B0(n25528), .B1(n28577), .Y(
        n24987) );
  AOI22XL U29683 ( .A0(n16659), .A1(n25526), .B0(n26262), .B1(n25532), .Y(
        n24984) );
  OAI211XL U29684 ( .A0(n25529), .A1(n16721), .B0(n24985), .C0(n24984), .Y(
        n24986) );
  NOR3XL U29685 ( .A(n24988), .B(n24987), .C(n24986), .Y(n25024) );
  OAI22XL U29686 ( .A0(n25140), .A1(n26274), .B0(n25522), .B1(n26279), .Y(
        n24993) );
  OAI22XL U29687 ( .A0(n25518), .A1(n28575), .B0(n25514), .B1(n28479), .Y(
        n24992) );
  OAI22XL U29688 ( .A0(n25513), .A1(n28577), .B0(n25515), .B1(n26285), .Y(
        n24991) );
  AOI22XL U29689 ( .A0(n36244), .A1(n25519), .B0(n26276), .B1(n25139), .Y(
        n24989) );
  OAI21XL U29690 ( .A0(n25141), .A1(n34958), .B0(n24989), .Y(n24990) );
  NOR4XL U29691 ( .A(n24993), .B(n24992), .C(n24991), .D(n24990), .Y(n25023)
         );
  OAI22XL U29692 ( .A0(n25543), .A1(n16661), .B0(n25541), .B1(n26274), .Y(
        n24998) );
  OAI2BB2XL U29693 ( .B0(n25163), .B1(n26285), .A0N(n25546), .A1N(n26262), .Y(
        n24997) );
  OAI22XL U29694 ( .A0(n25550), .A1(n28479), .B0(n25540), .B1(n28575), .Y(
        n24996) );
  AOI22XL U29695 ( .A0(n36244), .A1(n25542), .B0(n26276), .B1(n25545), .Y(
        n24994) );
  OAI2BB1XL U29696 ( .A0N(n16667), .A1N(n25547), .B0(n24994), .Y(n24995) );
  NOR4XL U29697 ( .A(n24998), .B(n24997), .C(n24996), .D(n24995), .Y(n25022)
         );
  OAI22XL U29698 ( .A0(n25587), .A1(n16661), .B0(n25586), .B1(n16721), .Y(
        n25003) );
  OAI22XL U29699 ( .A0(n25589), .A1(n26285), .B0(n25590), .B1(n28575), .Y(
        n25002) );
  AOI22XL U29700 ( .A0(n16659), .A1(n25588), .B0(n26276), .B1(n25585), .Y(
        n25000) );
  AOI22XL U29701 ( .A0(n26376), .A1(n25183), .B0(n26262), .B1(n25584), .Y(
        n24999) );
  OAI211XL U29702 ( .A0(n25597), .A1(n28577), .B0(n25000), .C0(n24999), .Y(
        n25001) );
  NOR3XL U29703 ( .A(n25003), .B(n25002), .C(n25001), .Y(n25054) );
  INVXL U29704 ( .A(n25004), .Y(n25605) );
  OAI22XL U29705 ( .A0(n25605), .A1(n26279), .B0(n25602), .B1(n16721), .Y(
        n25009) );
  OAI22XL U29706 ( .A0(n25603), .A1(n16661), .B0(n25604), .B1(n28575), .Y(
        n25008) );
  AOI22XL U29707 ( .A0(n16667), .A1(n25600), .B0(n26376), .B1(n25598), .Y(
        n25006) );
  AOI22XL U29708 ( .A0(n16659), .A1(n25601), .B0(n26276), .B1(n25599), .Y(
        n25005) );
  OAI211XL U29709 ( .A0(n25155), .A1(n26285), .B0(n25006), .C0(n25005), .Y(
        n25007) );
  NOR3XL U29710 ( .A(n25009), .B(n25008), .C(n25007), .Y(n25051) );
  AOI22XL U29711 ( .A0(n16667), .A1(n25563), .B0(n26376), .B1(n25010), .Y(
        n25016) );
  OAI22XL U29712 ( .A0(n25559), .A1(n26285), .B0(n25566), .B1(n16661), .Y(
        n25011) );
  AOI211XL U29713 ( .A0(n26262), .A1(n25561), .B0(n25012), .C0(n25011), .Y(
        n25014) );
  NAND2XL U29714 ( .A(n26276), .B(n25562), .Y(n25013) );
  NAND4XL U29715 ( .A(n25016), .B(n25015), .C(n25014), .D(n25013), .Y(n25052)
         );
  AOI22XL U29716 ( .A0(n36244), .A1(n25174), .B0(n16667), .B1(n25175), .Y(
        n25021) );
  OAI22XL U29717 ( .A0(n25575), .A1(n28575), .B0(n25574), .B1(n26285), .Y(
        n25019) );
  OAI22XL U29718 ( .A0(n25583), .A1(n28479), .B0(n25576), .B1(n26162), .Y(
        n25018) );
  OAI22XL U29719 ( .A0(n25573), .A1(n26274), .B0(n25177), .B1(n26279), .Y(
        n25017) );
  NOR3XL U29720 ( .A(n25019), .B(n25018), .C(n25017), .Y(n25020) );
  OAI211XL U29721 ( .A0(n25176), .A1(n34958), .B0(n25021), .C0(n25020), .Y(
        n25048) );
  NAND4XL U29722 ( .A(n25054), .B(n25051), .C(n25026), .D(n25025), .Y(n25027)
         );
  AOI2BB2XL U29723 ( .B0(n26276), .B1(n25621), .A0N(n28479), .A1N(n25623), .Y(
        n25035) );
  AOI22XL U29724 ( .A0(n28414), .A1(n25199), .B0(n26262), .B1(n25618), .Y(
        n25034) );
  OAI22XL U29725 ( .A0(n25620), .A1(n26274), .B0(n25622), .B1(n26285), .Y(
        n25032) );
  OAI22XL U29726 ( .A0(n25030), .A1(n28577), .B0(n16721), .B1(n25624), .Y(
        n25031) );
  AOI211XL U29727 ( .A0(n26263), .A1(n25628), .B0(n25032), .C0(n25031), .Y(
        n25033) );
  NAND3XL U29728 ( .A(n25035), .B(n25034), .C(n25033), .Y(n25057) );
  INVXL U29729 ( .A(n25205), .Y(n25633) );
  AOI22XL U29730 ( .A0(n16659), .A1(n25633), .B0(n26276), .B1(n25639), .Y(
        n25037) );
  AOI22XL U29731 ( .A0(n26263), .A1(n25632), .B0(n26262), .B1(n25638), .Y(
        n25036) );
  OAI211XL U29732 ( .A0(n25634), .A1(n26274), .B0(n25037), .C0(n25036), .Y(
        n25038) );
  AOI211XL U29733 ( .A0(n28556), .A1(n25635), .B0(n25039), .C0(n25038), .Y(
        n25041) );
  OAI211XL U29734 ( .A0(n25637), .A1(n26285), .B0(n25041), .C0(n25040), .Y(
        n25050) );
  OAI22XL U29735 ( .A0(n25653), .A1(n26162), .B0(n25652), .B1(n16721), .Y(
        n25045) );
  AOI22XL U29736 ( .A0(n16667), .A1(n25648), .B0(n26262), .B1(n25649), .Y(
        n25043) );
  NAND2XL U29737 ( .A(n26376), .B(n25647), .Y(n25042) );
  OAI211XL U29738 ( .A0(n25211), .A1(n26285), .B0(n25043), .C0(n25042), .Y(
        n25044) );
  NAND2XL U29739 ( .A(n28528), .B(n25657), .Y(n25046) );
  OAI211XL U29740 ( .A0(n25654), .A1(n34958), .B0(n25047), .C0(n25046), .Y(
        n25049) );
  NOR3XL U29741 ( .A(pool[49]), .B(n25050), .C(n25049), .Y(n25056) );
  NAND4BXL U29742 ( .AN(n25051), .B(n25050), .C(n25049), .D(n25048), .Y(n25053) );
  NAND4BBXL U29743 ( .AN(n25054), .BN(n25053), .C(pool[49]), .D(n25052), .Y(
        n25055) );
  NAND2XL U29744 ( .A(n34866), .B(pool[45]), .Y(n25060) );
  OAI21XL U29745 ( .A0(n25061), .A1(n34866), .B0(n25060), .Y(N29261) );
  OAI21XL U29746 ( .A0(conv_1[190]), .A1(n35363), .B0(n35365), .Y(n32989) );
  OAI2BB1XL U29747 ( .A0N(conv_1[190]), .A1N(n35364), .B0(n32988), .Y(n34085)
         );
  NAND2XL U29748 ( .A(n32989), .B(n34085), .Y(n25066) );
  NAND2XL U29749 ( .A(n32990), .B(n25066), .Y(n25065) );
  OAI211XL U29750 ( .A0(n32990), .A1(n25066), .B0(n33778), .C0(n25065), .Y(
        n25067) );
  OAI211XL U29751 ( .A0(n35368), .A1(n32990), .B0(n16652), .C0(n25067), .Y(
        n16272) );
  AOI22XL U29752 ( .A0(n33563), .A1(n25070), .B0(affine_1[28]), .B1(n25069), 
        .Y(n25071) );
  NAND2XL U29753 ( .A(n25071), .B(n33412), .Y(n16493) );
  NAND2XL U29754 ( .A(n27429), .B(n33990), .Y(n25072) );
  OAI21XL U29755 ( .A0(n33403), .A1(n33988), .B0(n25075), .Y(n27030) );
  INVXL U29756 ( .A(n25076), .Y(n25077) );
  NAND2XL U29757 ( .A(n35282), .B(conv_1[36]), .Y(n35288) );
  INVXL U29758 ( .A(conv_1[37]), .Y(n35291) );
  NAND2XL U29759 ( .A(n27301), .B(conv_1[38]), .Y(n27307) );
  OAI2BB1XL U29760 ( .A0N(n35295), .A1N(conv_1[40]), .B0(n35289), .Y(n35303)
         );
  OAI21XL U29761 ( .A0(conv_1[40]), .A1(n35294), .B0(n35296), .Y(n35301) );
  AOI22XL U29762 ( .A0(n32656), .A1(n25081), .B0(conv_1[42]), .B1(n25080), .Y(
        n25082) );
  NAND2XL U29763 ( .A(n25082), .B(n34682), .Y(n16421) );
  NOR4XL U29764 ( .A(in_data[8]), .B(in_data[7]), .C(in_data[13]), .D(
        in_data[9]), .Y(n25089) );
  OAI21XL U29765 ( .A0(in_data[1]), .A1(in_data[0]), .B0(in_data[2]), .Y(
        n25084) );
  NAND2XL U29766 ( .A(n25084), .B(n25083), .Y(n25086) );
  OR4XL U29767 ( .A(in_data[10]), .B(in_data[11]), .C(in_data[12]), .D(
        in_data[14]), .Y(n25085) );
  AOI31XL U29768 ( .A0(in_data[6]), .A1(in_data[5]), .A2(n25086), .B0(n25085), 
        .Y(n25088) );
  AOI32XL U29769 ( .A0(n25089), .A1(n22896), .A2(n25088), .B0(n25087), .B1(
        n23672), .Y(N17557) );
  INVXL U29770 ( .A(conv_1[113]), .Y(n25096) );
  NAND2XL U29771 ( .A(n34557), .B(n31343), .Y(n25092) );
  OAI21XL U29772 ( .A0(n34557), .A1(n31343), .B0(n25092), .Y(n25094) );
  AOI211XL U29773 ( .A0(n25096), .A1(n25094), .B0(n36042), .C0(n25093), .Y(
        n25095) );
  AOI2BB1XL U29774 ( .A0N(n25096), .A1N(n35330), .B0(n25095), .Y(n25097) );
  NAND2XL U29775 ( .A(n25097), .B(n34696), .Y(n16350) );
  AOI22XL U29776 ( .A0(n22362), .A1(n25098), .B0(n21100), .B1(n34929), .Y(
        n25099) );
  NAND2XL U29777 ( .A(n16721), .B(n34931), .Y(n25101) );
  NAND2XL U29778 ( .A(n25099), .B(n25101), .Y(n25461) );
  AOI22XL U29779 ( .A0(n22362), .A1(n34930), .B0(n21100), .B1(n25100), .Y(
        n25102) );
  NAND2XL U29780 ( .A(n25102), .B(n25101), .Y(n25460) );
  AOI222XL U29781 ( .A0(n25103), .A1(n28467), .B0(n25461), .B1(n28465), .C0(
        n25460), .C1(n35130), .Y(n25230) );
  AOI22XL U29782 ( .A0(n22362), .A1(n25105), .B0(n28407), .B1(n25104), .Y(
        n25106) );
  NAND2XL U29783 ( .A(n25106), .B(n25109), .Y(n25472) );
  AOI22XL U29784 ( .A0(n22362), .A1(n25108), .B0(n28407), .B1(n25107), .Y(
        n25110) );
  NAND2XL U29785 ( .A(n25110), .B(n25109), .Y(n25471) );
  AOI222XL U29786 ( .A0(n25111), .A1(n28467), .B0(n25472), .B1(n28465), .C0(
        n25471), .C1(n35130), .Y(n26350) );
  AOI22XL U29787 ( .A0(n22362), .A1(n25113), .B0(n25112), .B1(n25123), .Y(
        n25480) );
  AOI22XL U29788 ( .A0(n22362), .A1(n25115), .B0(n21100), .B1(n25114), .Y(
        n25117) );
  INVXL U29789 ( .A(n25116), .Y(n25484) );
  AOI222XL U29790 ( .A0(n25118), .A1(n28467), .B0(n35130), .B1(n25480), .C0(
        n25481), .C1(n16700), .Y(n34893) );
  AOI222XL U29791 ( .A0(n25230), .A1(pool[71]), .B0(n25230), .B1(n34893), .C0(
        pool[71]), .C1(n34893), .Y(n25129) );
  INVXL U29792 ( .A(pool[72]), .Y(n34895) );
  AOI211XL U29793 ( .A0(n28407), .A1(n25122), .B0(n25125), .C0(n25121), .Y(
        n25492) );
  OAI222XL U29794 ( .A0(n35135), .A1(n25492), .B0(n34989), .B1(n25493), .C0(
        n25128), .C1(N18471), .Y(n34894) );
  AOI222XL U29795 ( .A0(n25129), .A1(n34895), .B0(n25129), .B1(n34894), .C0(
        n34895), .C1(n34894), .Y(n25130) );
  AOI222XL U29796 ( .A0(n26350), .A1(pool[73]), .B0(n26350), .B1(n25130), .C0(
        pool[73]), .C1(n25130), .Y(n25198) );
  AOI22XL U29797 ( .A0(n22362), .A1(n25132), .B0(n21100), .B1(n25131), .Y(
        n25133) );
  NAND2XL U29798 ( .A(n25133), .B(n25136), .Y(n25506) );
  AOI22XL U29799 ( .A0(n22362), .A1(n25135), .B0(n21100), .B1(n25134), .Y(
        n25137) );
  NAND2XL U29800 ( .A(n25137), .B(n25136), .Y(n25505) );
  AOI222XL U29801 ( .A0(n25138), .A1(n28467), .B0(n25506), .B1(n28465), .C0(
        n25505), .C1(n35130), .Y(n26348) );
  AOI22XL U29802 ( .A0(n28528), .A1(n25139), .B0(n28571), .B1(n25519), .Y(
        n25146) );
  OAI22XL U29803 ( .A0(n25140), .A1(n16661), .B0(n25518), .B1(n35198), .Y(
        n25144) );
  OAI22XL U29804 ( .A0(n25141), .A1(n28553), .B0(n25513), .B1(n26621), .Y(
        n25143) );
  OAI22XL U29805 ( .A0(n25522), .A1(n28577), .B0(n25515), .B1(n34981), .Y(
        n25142) );
  NOR3XL U29806 ( .A(n25144), .B(n25143), .C(n25142), .Y(n25145) );
  OAI211XL U29807 ( .A0(n25514), .A1(n16672), .B0(n25146), .C0(n25145), .Y(
        n25194) );
  AOI22XL U29808 ( .A0(n28528), .A1(n25533), .B0(n28571), .B1(n25147), .Y(
        n25153) );
  AOI22XL U29809 ( .A0(n16660), .A1(n25531), .B0(n28559), .B1(n25526), .Y(
        n25152) );
  OAI22XL U29810 ( .A0(n25527), .A1(n28575), .B0(n25536), .B1(n16661), .Y(
        n25150) );
  OAI22XL U29811 ( .A0(n25148), .A1(n28553), .B0(n25528), .B1(n26621), .Y(
        n25149) );
  AOI211XL U29812 ( .A0(n28556), .A1(n25532), .B0(n25150), .C0(n25149), .Y(
        n25151) );
  NAND3XL U29813 ( .A(n25153), .B(n25152), .C(n25151), .Y(n25193) );
  OAI22XL U29814 ( .A0(n25605), .A1(n28577), .B0(n25154), .B1(n34958), .Y(
        n25161) );
  OAI22XL U29815 ( .A0(n25603), .A1(n28553), .B0(n25155), .B1(n34981), .Y(
        n25160) );
  AOI22XL U29816 ( .A0(n28528), .A1(n25599), .B0(n28559), .B1(n25601), .Y(
        n25158) );
  AOI22XL U29817 ( .A0(n28366), .A1(n25600), .B0(n28571), .B1(n25156), .Y(
        n25157) );
  OAI211XL U29818 ( .A0(n25604), .A1(n35198), .B0(n25158), .C0(n25157), .Y(
        n25159) );
  NOR3XL U29819 ( .A(n25161), .B(n25160), .C(n25159), .Y(n25220) );
  AOI22XL U29820 ( .A0(n16667), .A1(n25546), .B0(n18463), .B1(n25162), .Y(
        n25168) );
  AOI22XL U29821 ( .A0(n28324), .A1(n25547), .B0(n28571), .B1(n25542), .Y(
        n25167) );
  OAI22XL U29822 ( .A0(n25163), .A1(n28575), .B0(n25543), .B1(n28553), .Y(
        n25165) );
  OAI22XL U29823 ( .A0(n25541), .A1(n16661), .B0(n25540), .B1(n35198), .Y(
        n25164) );
  AOI211XL U29824 ( .A0(n34992), .A1(n25545), .B0(n25165), .C0(n25164), .Y(
        n25166) );
  NAND3XL U29825 ( .A(n25168), .B(n25167), .C(n25166), .Y(n25192) );
  AOI22XL U29826 ( .A0(n16660), .A1(n25558), .B0(n28571), .B1(n25560), .Y(
        n25173) );
  AOI22XL U29827 ( .A0(n28528), .A1(n25562), .B0(n28556), .B1(n25561), .Y(
        n25172) );
  OAI22XL U29828 ( .A0(n25559), .A1(n28575), .B0(n25566), .B1(n28553), .Y(
        n25170) );
  OAI22XL U29829 ( .A0(n25557), .A1(n34958), .B0(n25556), .B1(n16672), .Y(
        n25169) );
  AOI211XL U29830 ( .A0(n28324), .A1(n25563), .B0(n25170), .C0(n25169), .Y(
        n25171) );
  NAND3XL U29831 ( .A(n25173), .B(n25172), .C(n25171), .Y(n25221) );
  AOI22XL U29832 ( .A0(n28324), .A1(n25175), .B0(n28571), .B1(n25174), .Y(
        n25182) );
  OAI22XL U29833 ( .A0(n25573), .A1(n34958), .B0(n25176), .B1(n28553), .Y(
        n25180) );
  OAI22XL U29834 ( .A0(n25177), .A1(n28577), .B0(n25575), .B1(n35198), .Y(
        n25179) );
  OAI22XL U29835 ( .A0(n25574), .A1(n28575), .B0(n25583), .B1(n16672), .Y(
        n25178) );
  NOR3XL U29836 ( .A(n25180), .B(n25179), .C(n25178), .Y(n25181) );
  OAI211XL U29837 ( .A0(n25576), .A1(n28479), .B0(n25182), .C0(n25181), .Y(
        n25219) );
  AOI22XL U29838 ( .A0(n28528), .A1(n25585), .B0(n28559), .B1(n25588), .Y(
        n25189) );
  AOI22XL U29839 ( .A0(n26263), .A1(n25183), .B0(n16667), .B1(n25584), .Y(
        n25188) );
  OAI22XL U29840 ( .A0(n25589), .A1(n28575), .B0(n25597), .B1(n26621), .Y(
        n25185) );
  OAI22XL U29841 ( .A0(n28551), .A1(n25586), .B0(n25587), .B1(n28553), .Y(
        n25184) );
  AOI211XL U29842 ( .A0(n16660), .A1(n25186), .B0(n25185), .C0(n25184), .Y(
        n25187) );
  NAND3XL U29843 ( .A(n25189), .B(n25188), .C(n25187), .Y(n25218) );
  NOR4XL U29844 ( .A(n25192), .B(n25221), .C(n25219), .D(n25218), .Y(n25190)
         );
  NAND4XL U29845 ( .A(n26348), .B(n25191), .C(n25220), .D(n25190), .Y(n25197)
         );
  INVXL U29846 ( .A(n26348), .Y(n25195) );
  AOI22XL U29847 ( .A0(n28528), .A1(n25621), .B0(n28366), .B1(n25619), .Y(
        n25204) );
  AOI22XL U29848 ( .A0(n16660), .A1(n25199), .B0(n16670), .B1(n25628), .Y(
        n25203) );
  OAI22XL U29849 ( .A0(n28551), .A1(n25624), .B0(n25620), .B1(n16661), .Y(
        n25201) );
  OAI22XL U29850 ( .A0(n25623), .A1(n16672), .B0(n25622), .B1(n34981), .Y(
        n25200) );
  AOI211XL U29851 ( .A0(n28556), .A1(n25618), .B0(n25201), .C0(n25200), .Y(
        n25202) );
  NAND3XL U29852 ( .A(n25204), .B(n25203), .C(n25202), .Y(n25226) );
  AOI22XL U29853 ( .A0(n16660), .A1(n25643), .B0(n16670), .B1(n25632), .Y(
        n25210) );
  AOI22XL U29854 ( .A0(n28528), .A1(n25639), .B0(n28324), .B1(n25635), .Y(
        n25209) );
  OAI22XL U29855 ( .A0(n25637), .A1(n28575), .B0(n25634), .B1(n16661), .Y(
        n25207) );
  OAI22XL U29856 ( .A0(n28551), .A1(n25636), .B0(n25205), .B1(n16672), .Y(
        n25206) );
  AOI211XL U29857 ( .A0(n28556), .A1(n25638), .B0(n25207), .C0(n25206), .Y(
        n25208) );
  NAND3XL U29858 ( .A(n25210), .B(n25209), .C(n25208), .Y(n25217) );
  AOI22XL U29859 ( .A0(n26263), .A1(n25647), .B0(n16667), .B1(n25649), .Y(
        n25216) );
  AOI22XL U29860 ( .A0(n16660), .A1(n25651), .B0(n28559), .B1(n25657), .Y(
        n25215) );
  OAI22XL U29861 ( .A0(n25211), .A1(n28575), .B0(n25654), .B1(n28553), .Y(
        n25213) );
  OAI22XL U29862 ( .A0(n28551), .A1(n25652), .B0(n25653), .B1(n28479), .Y(
        n25212) );
  AOI211XL U29863 ( .A0(n28366), .A1(n25648), .B0(n25213), .C0(n25212), .Y(
        n25214) );
  NAND3XL U29864 ( .A(n25216), .B(n25215), .C(n25214), .Y(n25222) );
  NOR3XL U29865 ( .A(pool[74]), .B(n25217), .C(n25222), .Y(n25225) );
  NAND4BXL U29866 ( .AN(n25220), .B(n25219), .C(n25218), .D(n25217), .Y(n25223) );
  NAND4BXL U29867 ( .AN(n25223), .B(pool[74]), .C(n25222), .D(n25221), .Y(
        n25224) );
  NAND2XL U29868 ( .A(n34896), .B(pool[70]), .Y(n25229) );
  OAI21XL U29869 ( .A0(n25230), .A1(n34896), .B0(n25229), .Y(N29286) );
  NAND2BXL U29870 ( .AN(n25232), .B(n25231), .Y(n25234) );
  AOI211XL U29871 ( .A0(n25236), .A1(n25234), .B0(n36042), .C0(n25233), .Y(
        n25235) );
  AOI2BB1XL U29872 ( .A0N(n25236), .A1N(n35520), .B0(n25235), .Y(n25237) );
  NAND2XL U29873 ( .A(n25237), .B(n34689), .Y(n16021) );
  INVXL U29874 ( .A(conv_1[505]), .Y(n27130) );
  OAI31XL U29875 ( .A0(conv_1[503]), .A1(conv_1[504]), .A2(n27119), .B0(n27131), .Y(n27125) );
  OAI2BB1XL U29876 ( .A0N(n27130), .A1N(n27125), .B0(n27131), .Y(n27112) );
  NAND2XL U29877 ( .A(conv_1[503]), .B(n27119), .Y(n27118) );
  INVXL U29878 ( .A(n27131), .Y(n27120) );
  OAI2BB1XL U29879 ( .A0N(conv_1[505]), .A1N(n27126), .B0(n27120), .Y(n27132)
         );
  NAND2XL U29880 ( .A(n27112), .B(n27132), .Y(n25239) );
  AOI211XL U29881 ( .A0(n27113), .A1(n25239), .B0(n36042), .C0(n25238), .Y(
        n25240) );
  AOI2BB1XL U29882 ( .A0N(n27113), .A1N(n33427), .B0(n25240), .Y(n25241) );
  NAND2XL U29883 ( .A(n25241), .B(n34544), .Y(n15957) );
  AOI22XL U29884 ( .A0(n33563), .A1(n25244), .B0(affine_1[18]), .B1(n25243), 
        .Y(n25245) );
  NAND2XL U29885 ( .A(n25245), .B(n33564), .Y(n16483) );
  INVXL U29886 ( .A(conv_1[410]), .Y(n26520) );
  INVXL U29887 ( .A(conv_1[419]), .Y(n34675) );
  NAND4XL U29888 ( .A(conv_1[405]), .B(n27429), .C(n30672), .D(n34229), .Y(
        n25249) );
  NAND2XL U29889 ( .A(conv_1[405]), .B(n30672), .Y(n25248) );
  INVXL U29890 ( .A(n25248), .Y(n33520) );
  AOI221XL U29891 ( .A0(n35272), .A1(n25248), .B0(n27429), .B1(n33520), .C0(
        n28070), .Y(n31053) );
  NAND2XL U29892 ( .A(n31053), .B(conv_1[406]), .Y(n31052) );
  NAND2XL U29893 ( .A(n25249), .B(n31052), .Y(n30735) );
  AOI222XL U29894 ( .A0(n30736), .A1(conv_1[407]), .B0(n30736), .B1(n30735), 
        .C0(conv_1[407]), .C1(n30735), .Y(n25250) );
  INVXL U29895 ( .A(n25250), .Y(n25251) );
  NAND2XL U29896 ( .A(n34775), .B(n25253), .Y(n26521) );
  NAND2XL U29897 ( .A(n26521), .B(n26519), .Y(n25255) );
  AOI211XL U29898 ( .A0(n26520), .A1(n25255), .B0(n36042), .C0(n25254), .Y(
        n25256) );
  AOI2BB1XL U29899 ( .A0N(n26520), .A1N(n35487), .B0(n25256), .Y(n25257) );
  NAND2XL U29900 ( .A(n25257), .B(n34689), .Y(n16053) );
  INVXL U29901 ( .A(conv_1[522]), .Y(n29245) );
  INVXL U29902 ( .A(conv_1[520]), .Y(n30271) );
  NAND2XL U29903 ( .A(n25258), .B(conv_1[517]), .Y(n25261) );
  INVXL U29904 ( .A(conv_1[518]), .Y(n27259) );
  OAI21XL U29905 ( .A0(n30271), .A1(n30266), .B0(n30267), .Y(n35550) );
  AOI21XL U29906 ( .A0(n25262), .A1(n30266), .B0(n30267), .Y(n30265) );
  OAI21XL U29907 ( .A0(conv_1[520]), .A1(n30265), .B0(n29246), .Y(n35548) );
  NOR2BX1 U29908 ( .AN(n35548), .B(conv_1[521]), .Y(n35551) );
  AOI32XL U29909 ( .A0(conv_1[521]), .A1(n30267), .A2(n35550), .B0(n29246), 
        .B1(n35551), .Y(n25264) );
  AOI211XL U29910 ( .A0(n29245), .A1(n25264), .B0(n36042), .C0(n25263), .Y(
        n25265) );
  AOI2BB1XL U29911 ( .A0N(n29245), .A1N(n35547), .B0(n25265), .Y(n25266) );
  NAND2XL U29912 ( .A(n25266), .B(n34682), .Y(n15941) );
  NAND2XL U29913 ( .A(n34259), .B(n29383), .Y(n25267) );
  NAND2XL U29914 ( .A(n25270), .B(n25267), .Y(n25273) );
  INVXL U29915 ( .A(n25267), .Y(n25269) );
  AOI221XL U29916 ( .A0(n25274), .A1(n36020), .B0(n25269), .B1(n36020), .C0(
        n25268), .Y(n25271) );
  AOI2BB1XL U29917 ( .A0N(n25271), .A1N(n25270), .B0(n35549), .Y(n25272) );
  OAI31XL U29918 ( .A0(n25274), .A1(n36042), .A2(n25273), .B0(n25272), .Y(
        n16143) );
  NAND2XL U29919 ( .A(n25276), .B(n25275), .Y(n25278) );
  AOI211XL U29920 ( .A0(n25280), .A1(n25278), .B0(n36042), .C0(n25277), .Y(
        n25279) );
  AOI2BB1XL U29921 ( .A0N(n25280), .A1N(n35846), .B0(n25279), .Y(n25281) );
  NAND2XL U29922 ( .A(n25281), .B(n34408), .Y(n15235) );
  NAND2BXL U29923 ( .AN(n25283), .B(n25282), .Y(n25285) );
  AOI211XL U29924 ( .A0(n25287), .A1(n25285), .B0(n36042), .C0(n25284), .Y(
        n25286) );
  AOI2BB1XL U29925 ( .A0N(n25287), .A1N(n33863), .B0(n25286), .Y(n25288) );
  NAND2XL U29926 ( .A(n25288), .B(n34696), .Y(n16153) );
  AOI22XL U29927 ( .A0(n22762), .A1(conv_1[15]), .B0(n22690), .B1(conv_1[0]), 
        .Y(n25290) );
  NAND2XL U29928 ( .A(n25291), .B(n25290), .Y(n28406) );
  AOI22XL U29929 ( .A0(n22762), .A1(conv_1[135]), .B0(n16673), .B1(conv_1[165]), .Y(n25293) );
  AOI22XL U29930 ( .A0(n16662), .A1(conv_1[150]), .B0(n22616), .B1(conv_1[120]), .Y(n25292) );
  NAND2XL U29931 ( .A(n25293), .B(n25292), .Y(n34848) );
  INVXL U29932 ( .A(n34848), .Y(n26531) );
  AOI222XL U29933 ( .A0(n25294), .A1(n36246), .B0(n22690), .B1(conv_1[180]), 
        .C0(n22762), .C1(conv_1[195]), .Y(n34851) );
  OAI22XL U29934 ( .A0(n26531), .A1(n28577), .B0(n34851), .B1(n16661), .Y(
        n25311) );
  AOI22XL U29935 ( .A0(n16662), .A1(conv_1[390]), .B0(n16673), .B1(conv_1[405]), .Y(n25295) );
  NAND2XL U29936 ( .A(n25296), .B(n25295), .Y(n34824) );
  AOI222XL U29937 ( .A0(n25297), .A1(n36246), .B0(n18658), .B1(conv_1[420]), 
        .C0(n21011), .C1(conv_1[435]), .Y(n34823) );
  AOI222XL U29938 ( .A0(n25298), .A1(n22765), .B0(n16673), .B1(conv_1[285]), 
        .C0(conv_1[270]), .C1(n25289), .Y(n34822) );
  AOI22XL U29939 ( .A0(n16662), .A1(conv_1[330]), .B0(n25299), .B1(conv_1[300]), .Y(n25300) );
  NAND2XL U29940 ( .A(n25301), .B(n25300), .Y(n34825) );
  OAI2BB2XL U29941 ( .B0(n34822), .B1(n25402), .A0N(n34825), .A1N(n28289), .Y(
        n25302) );
  AOI211XL U29942 ( .A0(n25399), .A1(n34824), .B0(n25303), .C0(n25302), .Y(
        n28404) );
  NAND2XL U29943 ( .A(n36244), .B(n34847), .Y(n28403) );
  AOI22XL U29944 ( .A0(n25299), .A1(conv_1[60]), .B0(n16673), .B1(conv_1[105]), 
        .Y(n25308) );
  NAND2XL U29945 ( .A(n25308), .B(n25307), .Y(n34846) );
  NAND2XL U29946 ( .A(n16659), .B(n34846), .Y(n25309) );
  OAI211XL U29947 ( .A0(n28404), .A1(n28467), .B0(n28403), .C0(n25309), .Y(
        n25310) );
  OAI22XL U29948 ( .A0(n28416), .A1(n26162), .B0(n28415), .B1(n26274), .Y(
        n25317) );
  AOI22XL U29949 ( .A0(n28556), .A1(n25312), .B0(n26262), .B1(n28411), .Y(
        n25315) );
  AOI22XL U29950 ( .A0(n36244), .A1(n28421), .B0(n28413), .B1(n26260), .Y(
        n25313) );
  NAND3XL U29951 ( .A(n25315), .B(n25314), .C(n25313), .Y(n25316) );
  AOI22XL U29952 ( .A0(n28528), .A1(n26586), .B0(n26276), .B1(n28499), .Y(
        n25322) );
  OAI22XL U29953 ( .A0(n28501), .A1(n26274), .B0(n28504), .B1(n26285), .Y(
        n25320) );
  INVXL U29954 ( .A(n28498), .Y(n26422) );
  OAI22XL U29955 ( .A0(n28502), .A1(n16661), .B0(n26422), .B1(n28577), .Y(
        n25319) );
  OAI22XL U29956 ( .A0(n28503), .A1(n28575), .B0(n28511), .B1(n16721), .Y(
        n25318) );
  NOR3XL U29957 ( .A(n25320), .B(n25319), .C(n25318), .Y(n25321) );
  OAI211XL U29958 ( .A0(n28500), .A1(n26279), .B0(n25322), .C0(n25321), .Y(
        n25370) );
  AOI22XL U29959 ( .A0(n36244), .A1(n26585), .B0(n16667), .B1(n28475), .Y(
        n25326) );
  OAI22XL U29960 ( .A0(n28472), .A1(n16661), .B0(n28471), .B1(n26285), .Y(
        n25324) );
  OAI22XL U29961 ( .A0(n28469), .A1(n26274), .B0(n28480), .B1(n26162), .Y(
        n25323) );
  AOI211XL U29962 ( .A0(n34992), .A1(n28473), .B0(n25324), .C0(n25323), .Y(
        n25325) );
  NAND3XL U29963 ( .A(n25327), .B(n25326), .C(n25325), .Y(n25369) );
  AOI22XL U29964 ( .A0(n26263), .A1(n26595), .B0(n26262), .B1(n28484), .Y(
        n25333) );
  AOI22XL U29965 ( .A0(n36244), .A1(n28494), .B0(n28528), .B1(n28486), .Y(
        n25332) );
  OAI22XL U29966 ( .A0(n28491), .A1(n28575), .B0(n28490), .B1(n26285), .Y(
        n25328) );
  AOI211XL U29967 ( .A0(n16667), .A1(n28487), .B0(n25329), .C0(n25328), .Y(
        n25331) );
  NAND2XL U29968 ( .A(n26276), .B(n28485), .Y(n25330) );
  NAND4XL U29969 ( .A(n25333), .B(n25332), .C(n25331), .D(n25330), .Y(n25358)
         );
  AOI22XL U29970 ( .A0(n16667), .A1(n26570), .B0(n26172), .B1(n26411), .Y(
        n25344) );
  AOI22XL U29971 ( .A0(n25337), .A1(n26413), .B0(n25336), .B1(n25335), .Y(
        n25341) );
  AOI22XL U29972 ( .A0(n25399), .A1(n25339), .B0(n28289), .B1(n25338), .Y(
        n25340) );
  OAI211XL U29973 ( .A0(n26410), .A1(n16721), .B0(n25341), .C0(n25340), .Y(
        n28468) );
  AOI22XL U29974 ( .A0(N18471), .A1(n28468), .B0(n28528), .B1(n26569), .Y(
        n25342) );
  NAND3XL U29975 ( .A(n25344), .B(n25343), .C(n25342), .Y(n34794) );
  NAND4XL U29976 ( .A(n25370), .B(n25369), .C(n25358), .D(n34794), .Y(n25411)
         );
  AOI22XL U29977 ( .A0(n26263), .A1(n28437), .B0(n26376), .B1(n25345), .Y(
        n25351) );
  OAI22XL U29978 ( .A0(n28443), .A1(n26162), .B0(n28442), .B1(n26279), .Y(
        n25349) );
  OAI22XL U29979 ( .A0(n28438), .A1(n28479), .B0(n28449), .B1(n28575), .Y(
        n25348) );
  OAI22XL U29980 ( .A0(n28439), .A1(n26285), .B0(n25346), .B1(n16721), .Y(
        n25347) );
  NOR3XL U29981 ( .A(n25349), .B(n25348), .C(n25347), .Y(n25350) );
  OAI211XL U29982 ( .A0(n28440), .A1(n28577), .B0(n25351), .C0(n25350), .Y(
        n25423) );
  AOI22XL U29983 ( .A0(n36244), .A1(n26609), .B0(n16667), .B1(n28514), .Y(
        n25353) );
  OAI211XL U29984 ( .A0(n28516), .A1(n26274), .B0(n25353), .C0(n25352), .Y(
        n25354) );
  AOI211XL U29985 ( .A0(n34992), .A1(n28512), .B0(n25355), .C0(n25354), .Y(
        n25357) );
  NAND2XL U29986 ( .A(n26276), .B(n28522), .Y(n25356) );
  OAI211XL U29987 ( .A0(n28519), .A1(n34958), .B0(n25357), .C0(n25356), .Y(
        n25429) );
  NOR4XL U29988 ( .A(n25423), .B(n25358), .C(n34794), .D(n25429), .Y(n25372)
         );
  INVXL U29989 ( .A(n28456), .Y(n26450) );
  AOI22XL U29990 ( .A0(n36244), .A1(n28450), .B0(n26263), .B1(n26450), .Y(
        n25363) );
  OAI22XL U29991 ( .A0(n28454), .A1(n26279), .B0(n28463), .B1(n28575), .Y(
        n25361) );
  OAI22XL U29992 ( .A0(n28452), .A1(n26162), .B0(n26452), .B1(n28577), .Y(
        n25360) );
  OAI22XL U29993 ( .A0(n28453), .A1(n26274), .B0(n28457), .B1(n28479), .Y(
        n25359) );
  NOR3XL U29994 ( .A(n25361), .B(n25360), .C(n25359), .Y(n25362) );
  OAI211XL U29995 ( .A0(n28455), .A1(n26285), .B0(n25363), .C0(n25362), .Y(
        n25424) );
  AOI22XL U29996 ( .A0(n28528), .A1(n28529), .B0(n16667), .B1(n28530), .Y(
        n25368) );
  OAI22XL U29997 ( .A0(n28531), .A1(n26274), .B0(n28534), .B1(n16721), .Y(
        n25365) );
  OAI22XL U29998 ( .A0(n28532), .A1(n26285), .B0(n28533), .B1(n34958), .Y(
        n25364) );
  AOI211XL U29999 ( .A0(n26262), .A1(n28537), .B0(n25365), .C0(n25364), .Y(
        n25366) );
  NAND3XL U30000 ( .A(n25368), .B(n25367), .C(n25366), .Y(n25425) );
  NOR4XL U30001 ( .A(n25370), .B(n25424), .C(n25369), .D(n25425), .Y(n25371)
         );
  AOI21XL U30002 ( .A0(n25372), .A1(n25371), .B0(pool[4]), .Y(n25410) );
  OAI22XL U30003 ( .A0(n25376), .A1(n25402), .B0(n25375), .B1(n25393), .Y(
        n25377) );
  AOI22XL U30004 ( .A0(N18471), .A1(n28427), .B0(n16667), .B1(n26538), .Y(
        n25381) );
  NAND2XL U30005 ( .A(n25382), .B(n25381), .Y(n25383) );
  INVXL U30006 ( .A(n26563), .Y(n26400) );
  NAND2XL U30007 ( .A(n36244), .B(n26562), .Y(n25390) );
  OAI2BB1XL U30008 ( .A0N(n28289), .A1N(n25384), .B0(n25390), .Y(n25386) );
  OAI22XL U30009 ( .A0(n26566), .A1(n25402), .B0(n26401), .B1(n25393), .Y(
        n25385) );
  OAI22XL U30010 ( .A0(n28428), .A1(n28467), .B0(n26556), .B1(n28479), .Y(
        n25388) );
  NAND2XL U30011 ( .A(n25400), .B(n26172), .Y(n26390) );
  INVXL U30012 ( .A(n26390), .Y(n25406) );
  OAI22XL U30013 ( .A0(n25396), .A1(n25395), .B0(n25394), .B1(n25393), .Y(
        n25397) );
  NAND2XL U30014 ( .A(n36244), .B(n25400), .Y(n26392) );
  OAI211XL U30015 ( .A0(n26393), .A1(n25402), .B0(n25401), .C0(n26392), .Y(
        n28433) );
  AOI22XL U30016 ( .A0(N18471), .A1(n28433), .B0(n16667), .B1(n26547), .Y(
        n25403) );
  NAND2XL U30017 ( .A(n25404), .B(n25403), .Y(n25405) );
  AOI222XL U30018 ( .A0(pool[0]), .A1(pool[1]), .B0(pool[0]), .B1(n34790), 
        .C0(pool[1]), .C1(n34790), .Y(n25407) );
  AOI222XL U30019 ( .A0(n34793), .A1(n34792), .B0(n34793), .B1(n25407), .C0(
        n34792), .C1(n25407), .Y(n25408) );
  AOI222XL U30020 ( .A0(n25685), .A1(pool[3]), .B0(n25685), .B1(n25408), .C0(
        pool[3]), .C1(n25408), .Y(n25409) );
  OAI22XL U30021 ( .A0(n28550), .A1(n16721), .B0(n28552), .B1(n28575), .Y(
        n25416) );
  OAI22XL U30022 ( .A0(n28554), .A1(n16661), .B0(n28563), .B1(n26285), .Y(
        n25415) );
  AOI22XL U30023 ( .A0(n34992), .A1(n28558), .B0(n26262), .B1(n28555), .Y(
        n25413) );
  AOI22XL U30024 ( .A0(n16667), .A1(n28560), .B0(n26276), .B1(n28557), .Y(
        n25412) );
  OAI211XL U30025 ( .A0(n28549), .A1(n26274), .B0(n25413), .C0(n25412), .Y(
        n25414) );
  NOR3XL U30026 ( .A(n25416), .B(n25415), .C(n25414), .Y(n25428) );
  OAI22XL U30027 ( .A0(n28576), .A1(n26285), .B0(n28580), .B1(n26274), .Y(
        n25422) );
  OAI22XL U30028 ( .A0(n26642), .A1(n16721), .B0(n28579), .B1(n28479), .Y(
        n25421) );
  OAI22XL U30029 ( .A0(n28578), .A1(n26279), .B0(n25417), .B1(n34958), .Y(
        n25420) );
  AOI22XL U30030 ( .A0(n16667), .A1(n28573), .B0(n26276), .B1(n28572), .Y(
        n25418) );
  OAI2BB1X1 U30031 ( .A0N(n34963), .A1N(n28574), .B0(n25418), .Y(n25419) );
  NAND3XL U30032 ( .A(n25428), .B(n25427), .C(n34796), .Y(n25431) );
  NAND4XL U30033 ( .A(pool[4]), .B(n25425), .C(n25424), .D(n25423), .Y(n25426)
         );
  NAND2XL U30034 ( .A(n34795), .B(pool[0]), .Y(n25435) );
  OAI21XL U30035 ( .A0(n25436), .A1(n34795), .B0(n25435), .Y(N29216) );
  AOI21XL U30036 ( .A0(conv_1[220]), .A1(n25438), .B0(n35392), .Y(n28600) );
  OAI21XL U30037 ( .A0(n25440), .A1(n16655), .B0(n35395), .Y(n25439) );
  NAND2XL U30038 ( .A(n25442), .B(n34544), .Y(n16242) );
  AOI22XL U30039 ( .A0(n34864), .A1(n25444), .B0(n25443), .B1(n34866), .Y(
        N29265) );
  AOI22XL U30040 ( .A0(n34864), .A1(n25446), .B0(n25445), .B1(n34866), .Y(
        N29264) );
  INVXL U30041 ( .A(conv_1[131]), .Y(n25452) );
  NAND2XL U30042 ( .A(n34292), .B(n30450), .Y(n25448) );
  OAI21XL U30043 ( .A0(n34292), .A1(n30450), .B0(n25448), .Y(n25450) );
  AOI211XL U30044 ( .A0(n25452), .A1(n25450), .B0(n36042), .C0(n25449), .Y(
        n25451) );
  AOI2BB1XL U30045 ( .A0N(n25452), .A1N(n34296), .B0(n25451), .Y(n25453) );
  NAND2XL U30046 ( .A(n25453), .B(n34682), .Y(n16332) );
  AOI32XL U30047 ( .A0(n34461), .A1(n35676), .A2(n25454), .B0(n16655), .B1(
        n35676), .Y(n25455) );
  AOI32XL U30048 ( .A0(n34461), .A1(n25456), .A2(n34742), .B0(conv_3[225]), 
        .B1(n25455), .Y(n25457) );
  NAND2XL U30049 ( .A(n25457), .B(n34755), .Y(n15908) );
  OAI22XL U30050 ( .A0(n25459), .A1(n35200), .B0(n25458), .B1(n28349), .Y(
        n25466) );
  AOI22XL U30051 ( .A0(n25766), .A1(n34931), .B0(n28366), .B1(n34932), .Y(
        n25463) );
  AOI22XL U30052 ( .A0(n35130), .A1(n25461), .B0(n34827), .B1(n25460), .Y(
        n25462) );
  OAI211XL U30053 ( .A0(n25464), .A1(n28553), .B0(n25463), .C0(n25462), .Y(
        n25465) );
  AOI22XL U30054 ( .A0(n16665), .A1(n25468), .B0(n16664), .B1(n25467), .Y(
        n25476) );
  AOI22XL U30055 ( .A0(n28366), .A1(n25470), .B0(n16663), .B1(n25469), .Y(
        n25475) );
  AOI22XL U30056 ( .A0(n35130), .A1(n25472), .B0(n34827), .B1(n25471), .Y(
        n25474) );
  AOI22XL U30057 ( .A0(n16665), .A1(n25479), .B0(n16664), .B1(n25478), .Y(
        n25483) );
  AOI22XL U30058 ( .A0(n35130), .A1(n25481), .B0(n34827), .B1(n25480), .Y(
        n25482) );
  OAI211XL U30059 ( .A0(n35135), .A1(n25484), .B0(n25483), .C0(n25482), .Y(
        n25485) );
  AOI222XL U30060 ( .A0(n25674), .A1(pool[76]), .B0(n25674), .B1(n34898), .C0(
        pool[76]), .C1(n34898), .Y(n25499) );
  AOI22XL U30061 ( .A0(n16665), .A1(n25489), .B0(n16664), .B1(n25488), .Y(
        n25498) );
  OAI22XL U30062 ( .A0(n25491), .A1(n26621), .B0(n25490), .B1(n28349), .Y(
        n25495) );
  OAI22XL U30063 ( .A0(n25493), .A1(n26575), .B0(n25492), .B1(n34989), .Y(
        n25494) );
  AOI222XL U30064 ( .A0(n25499), .A1(n34899), .B0(n25499), .B1(n34900), .C0(
        n34899), .C1(n34900), .Y(n25500) );
  AOI222XL U30065 ( .A0(pool[78]), .A1(n27369), .B0(pool[78]), .B1(n25500), 
        .C0(n27369), .C1(n25500), .Y(n25617) );
  OAI2BB2XL U30066 ( .B0(n25502), .B1(n26621), .A0N(n25501), .A1N(n25766), .Y(
        n25510) );
  AOI22XL U30067 ( .A0(n16665), .A1(n25504), .B0(n16664), .B1(n25503), .Y(
        n25508) );
  AOI22XL U30068 ( .A0(n35130), .A1(n25506), .B0(n34827), .B1(n25505), .Y(
        n25507) );
  NAND2XL U30069 ( .A(n25508), .B(n25507), .Y(n25509) );
  AOI211XL U30070 ( .A0(n16663), .A1(n25511), .B0(n25510), .C0(n25509), .Y(
        n27371) );
  OAI22XL U30071 ( .A0(n25513), .A1(n35198), .B0(n25512), .B1(n28553), .Y(
        n25525) );
  OAI22XL U30072 ( .A0(n25515), .A1(n26621), .B0(n25514), .B1(n18208), .Y(
        n25524) );
  AOI22XL U30073 ( .A0(n28559), .A1(n25517), .B0(n16663), .B1(n25516), .Y(
        n25521) );
  AOI2BB2XL U30074 ( .B0(n25795), .B1(n25519), .A0N(n35239), .A1N(n25518), .Y(
        n25520) );
  OAI211XL U30075 ( .A0(n25522), .A1(n35200), .B0(n25521), .C0(n25520), .Y(
        n25523) );
  NOR3XL U30076 ( .A(n25525), .B(n25524), .C(n25523), .Y(n25555) );
  OAI2BB2XL U30077 ( .B0(n25527), .B1(n26621), .A0N(n25526), .A1N(n35236), .Y(
        n25539) );
  OAI22XL U30078 ( .A0(n25529), .A1(n25771), .B0(n25528), .B1(n35198), .Y(
        n25538) );
  AOI22XL U30079 ( .A0(n35195), .A1(n25531), .B0(n28559), .B1(n25530), .Y(
        n25535) );
  AOI22XL U30080 ( .A0(n16665), .A1(n25533), .B0(n16664), .B1(n25532), .Y(
        n25534) );
  OAI211XL U30081 ( .A0(n25536), .A1(n28349), .B0(n25535), .C0(n25534), .Y(
        n25537) );
  NOR3XL U30082 ( .A(n25539), .B(n25538), .C(n25537), .Y(n25554) );
  OAI22XL U30083 ( .A0(n25541), .A1(n28349), .B0(n25540), .B1(n35239), .Y(
        n25553) );
  OAI2BB2XL U30084 ( .B0(n25543), .B1(n16672), .A0N(n25542), .A1N(n25795), .Y(
        n25552) );
  AOI22XL U30085 ( .A0(n16665), .A1(n25545), .B0(n28366), .B1(n25544), .Y(
        n25549) );
  AOI22XL U30086 ( .A0(n16660), .A1(n25547), .B0(n16664), .B1(n25546), .Y(
        n25548) );
  OAI211XL U30087 ( .A0(n25550), .A1(n18208), .B0(n25549), .C0(n25548), .Y(
        n25551) );
  NOR3XL U30088 ( .A(n25553), .B(n25552), .C(n25551), .Y(n25612) );
  AND2XL U30089 ( .A(n25555), .B(n25554), .Y(n25614) );
  OAI22XL U30090 ( .A0(n25557), .A1(n28349), .B0(n25556), .B1(n18208), .Y(
        n25569) );
  OAI2BB2XL U30091 ( .B0(n25559), .B1(n26621), .A0N(n25558), .A1N(n35195), .Y(
        n25568) );
  AOI22XL U30092 ( .A0(n16664), .A1(n25561), .B0(n25795), .B1(n25560), .Y(
        n25565) );
  AOI22XL U30093 ( .A0(n16660), .A1(n25563), .B0(n16670), .B1(n25562), .Y(
        n25564) );
  OAI211XL U30094 ( .A0(n25566), .A1(n16672), .B0(n25565), .C0(n25564), .Y(
        n25567) );
  NOR3XL U30095 ( .A(n25569), .B(n25568), .C(n25567), .Y(n25664) );
  AOI22XL U30096 ( .A0(n28559), .A1(n25571), .B0(n16664), .B1(n25570), .Y(
        n25582) );
  OAI22XL U30097 ( .A0(n25573), .A1(n28349), .B0(n25572), .B1(n35198), .Y(
        n25580) );
  OAI22XL U30098 ( .A0(n25575), .A1(n35239), .B0(n25574), .B1(n26621), .Y(
        n25579) );
  OAI22XL U30099 ( .A0(n25577), .A1(n25771), .B0(n25576), .B1(n28553), .Y(
        n25578) );
  NOR3XL U30100 ( .A(n25580), .B(n25579), .C(n25578), .Y(n25581) );
  OAI211XL U30101 ( .A0(n25583), .A1(n18208), .B0(n25582), .C0(n25581), .Y(
        n25665) );
  AOI22XL U30102 ( .A0(n16665), .A1(n25585), .B0(n16664), .B1(n25584), .Y(
        n25596) );
  OAI22XL U30103 ( .A0(n25587), .A1(n16672), .B0(n25586), .B1(n25771), .Y(
        n25594) );
  OAI2BB2XL U30104 ( .B0(n25589), .B1(n26621), .A0N(n25588), .A1N(n35236), .Y(
        n25593) );
  OAI22XL U30105 ( .A0(n25591), .A1(n28349), .B0(n25590), .B1(n35239), .Y(
        n25592) );
  NOR3XL U30106 ( .A(n25594), .B(n25593), .C(n25592), .Y(n25595) );
  OAI211XL U30107 ( .A0(n25597), .A1(n35198), .B0(n25596), .C0(n25595), .Y(
        n25663) );
  AOI22XL U30108 ( .A0(n16665), .A1(n25599), .B0(n16663), .B1(n25598), .Y(
        n25611) );
  AOI22XL U30109 ( .A0(n35236), .A1(n25601), .B0(n16660), .B1(n25600), .Y(
        n25610) );
  OAI22XL U30110 ( .A0(n25603), .A1(n16672), .B0(n25602), .B1(n25771), .Y(
        n25607) );
  OAI22XL U30111 ( .A0(n25605), .A1(n35200), .B0(n25604), .B1(n35239), .Y(
        n25606) );
  AOI211XL U30112 ( .A0(n28324), .A1(n25608), .B0(n25607), .C0(n25606), .Y(
        n25609) );
  NAND3XL U30113 ( .A(n25611), .B(n25610), .C(n25609), .Y(n25662) );
  NOR4BXL U30114 ( .AN(n25612), .B(n25665), .C(n25663), .D(n25662), .Y(n25613)
         );
  NAND4XL U30115 ( .A(n27371), .B(n25614), .C(n25664), .D(n25613), .Y(n25615)
         );
  AOI22XL U30116 ( .A0(n16660), .A1(n25619), .B0(n16664), .B1(n25618), .Y(
        n25631) );
  AOI2BB2XL U30117 ( .B0(n16670), .B1(n25621), .A0N(n28349), .A1N(n25620), .Y(
        n25630) );
  OAI22XL U30118 ( .A0(n25623), .A1(n18208), .B0(n25622), .B1(n26621), .Y(
        n25627) );
  OAI22XL U30119 ( .A0(n25625), .A1(n35239), .B0(n25624), .B1(n25771), .Y(
        n25626) );
  AOI211XL U30120 ( .A0(n18463), .A1(n25628), .B0(n25627), .C0(n25626), .Y(
        n25629) );
  NAND3XL U30121 ( .A(n25631), .B(n25630), .C(n25629), .Y(n25670) );
  AOI22XL U30122 ( .A0(n35236), .A1(n25633), .B0(n18463), .B1(n25632), .Y(
        n25646) );
  AOI2BB2XL U30123 ( .B0(n16660), .B1(n25635), .A0N(n28349), .A1N(n25634), .Y(
        n25645) );
  OAI22XL U30124 ( .A0(n25637), .A1(n26621), .B0(n25636), .B1(n25771), .Y(
        n25642) );
  AOI22XL U30125 ( .A0(n25639), .A1(n16670), .B0(n25638), .B1(n16664), .Y(
        n25640) );
  INVXL U30126 ( .A(n25640), .Y(n25641) );
  AOI211XL U30127 ( .A0(n35195), .A1(n25643), .B0(n25642), .C0(n25641), .Y(
        n25644) );
  NAND3XL U30128 ( .A(n25646), .B(n25645), .C(n25644), .Y(n25661) );
  AOI22XL U30129 ( .A0(n16660), .A1(n25648), .B0(n16663), .B1(n25647), .Y(
        n25660) );
  AOI22XL U30130 ( .A0(n28324), .A1(n25650), .B0(n16664), .B1(n25649), .Y(
        n25659) );
  OAI2BB2XL U30131 ( .B0(n25652), .B1(n25771), .A0N(n25651), .A1N(n35195), .Y(
        n25656) );
  OAI22XL U30132 ( .A0(n25654), .A1(n16672), .B0(n25653), .B1(n28553), .Y(
        n25655) );
  AOI211XL U30133 ( .A0(n35236), .A1(n25657), .B0(n25656), .C0(n25655), .Y(
        n25658) );
  NAND3XL U30134 ( .A(n25660), .B(n25659), .C(n25658), .Y(n25666) );
  NOR3XL U30135 ( .A(pool[79]), .B(n25661), .C(n25666), .Y(n25669) );
  NAND4BXL U30136 ( .AN(n25664), .B(n25663), .C(n25662), .D(n25661), .Y(n25667) );
  NAND4BXL U30137 ( .AN(n25667), .B(pool[79]), .C(n25666), .D(n25665), .Y(
        n25668) );
  NAND2XL U30138 ( .A(n34901), .B(pool[75]), .Y(n25673) );
  OAI21XL U30139 ( .A0(n25674), .A1(n34901), .B0(n25673), .Y(N29291) );
  INVXL U30140 ( .A(conv_2[109]), .Y(n34407) );
  NAND2XL U30141 ( .A(n29046), .B(n34717), .Y(n25678) );
  AOI222XL U30142 ( .A0(n27139), .A1(n27140), .B0(n27139), .B1(conv_2[108]), 
        .C0(n27140), .C1(conv_2[108]), .Y(n25677) );
  NAND2XL U30143 ( .A(n25678), .B(n25677), .Y(n34403) );
  NAND2XL U30144 ( .A(n35884), .B(n25679), .Y(n28680) );
  NAND2XL U30145 ( .A(n28678), .B(n28680), .Y(n25681) );
  AOI211XL U30146 ( .A0(n28679), .A1(n25681), .B0(n16655), .C0(n25680), .Y(
        n25682) );
  AOI2BB1XL U30147 ( .A0N(n28679), .A1N(n35894), .B0(n25682), .Y(n25683) );
  NAND2XL U30148 ( .A(n25683), .B(n35859), .Y(n15133) );
  INVXL U30149 ( .A(n34795), .Y(n34791) );
  AOI22XL U30150 ( .A0(n34791), .A1(n25685), .B0(n25684), .B1(n34795), .Y(
        N29219) );
  OAI22XL U30151 ( .A0(n28288), .A1(n28349), .B0(n28285), .B1(n26621), .Y(
        n25690) );
  AOI22XL U30152 ( .A0(n25766), .A1(n35230), .B0(n16664), .B1(n28294), .Y(
        n25687) );
  NAND2XL U30153 ( .A(n16670), .B(n28293), .Y(n25686) );
  OAI211XL U30154 ( .A0(n25688), .A1(n16701), .B0(n25687), .C0(n25686), .Y(
        n25689) );
  AOI22XL U30155 ( .A0(n16664), .A1(n26166), .B0(n25795), .B1(n35169), .Y(
        n25696) );
  AOI22XL U30156 ( .A0(n35195), .A1(n28265), .B0(n18463), .B1(n35167), .Y(
        n25695) );
  OAI22XL U30157 ( .A0(n35170), .A1(n26621), .B0(n35172), .B1(n35198), .Y(
        n25693) );
  OAI22XL U30158 ( .A0(n26163), .A1(n28553), .B0(n35171), .B1(n28349), .Y(
        n25692) );
  AOI211XL U30159 ( .A0(n35236), .A1(n35168), .B0(n25693), .C0(n25692), .Y(
        n25694) );
  NAND3XL U30160 ( .A(n25696), .B(n25695), .C(n25694), .Y(n25808) );
  OAI22XL U30161 ( .A0(n25698), .A1(n26621), .B0(n25697), .B1(n28349), .Y(
        n25705) );
  AOI22XL U30162 ( .A0(n16665), .A1(n25700), .B0(n16664), .B1(n25699), .Y(
        n25702) );
  NAND2XL U30163 ( .A(n28465), .B(n25701), .Y(n28270) );
  OAI211XL U30164 ( .A0(n25703), .A1(n16701), .B0(n25702), .C0(n28270), .Y(
        n25704) );
  AOI22XL U30165 ( .A0(n25766), .A1(n35153), .B0(n16670), .B1(n25707), .Y(
        n25711) );
  AOI22XL U30166 ( .A0(n35130), .A1(n25709), .B0(n34827), .B1(n25708), .Y(
        n25710) );
  OAI211XL U30167 ( .A0(n25712), .A1(n28349), .B0(n25711), .C0(n25710), .Y(
        n25713) );
  AOI222XL U30168 ( .A0(n25811), .A1(pool[121]), .B0(n25811), .B1(n26702), 
        .C0(pool[121]), .C1(n26702), .Y(n25724) );
  AOI22XL U30169 ( .A0(n28366), .A1(n35139), .B0(n16663), .B1(n28279), .Y(
        n25723) );
  AOI22XL U30170 ( .A0(n16665), .A1(n25717), .B0(n16664), .B1(n25716), .Y(
        n25722) );
  AOI22XL U30171 ( .A0(n35130), .A1(n25719), .B0(n34827), .B1(n25718), .Y(
        n25721) );
  OR2XL U30172 ( .A(n35241), .B(n25720), .Y(n28275) );
  AOI222XL U30173 ( .A0(n25724), .A1(n35021), .B0(n25724), .B1(n35020), .C0(
        n35021), .C1(n35020), .Y(n25725) );
  AOI222XL U30174 ( .A0(n26704), .A1(pool[123]), .B0(n26704), .B1(n25725), 
        .C0(pool[123]), .C1(n25725), .Y(n25785) );
  AOI22XL U30175 ( .A0(n16663), .A1(n28352), .B0(n16664), .B1(n26237), .Y(
        n25731) );
  AOI22XL U30176 ( .A0(n16660), .A1(n28351), .B0(n16670), .B1(n26240), .Y(
        n25730) );
  OAI22XL U30177 ( .A0(n35053), .A1(n26621), .B0(n25726), .B1(n18208), .Y(
        n25728) );
  OAI22XL U30178 ( .A0(n35057), .A1(n16672), .B0(n35055), .B1(n35239), .Y(
        n25727) );
  AOI211XL U30179 ( .A0(n25795), .A1(n35054), .B0(n25728), .C0(n25727), .Y(
        n25729) );
  NAND3XL U30180 ( .A(n25731), .B(n25730), .C(n25729), .Y(n25794) );
  AOI22XL U30181 ( .A0(n16664), .A1(n26244), .B0(n25795), .B1(n35034), .Y(
        n25737) );
  AOI22XL U30182 ( .A0(n35236), .A1(n35040), .B0(n18197), .B1(n28344), .Y(
        n25736) );
  OAI22XL U30183 ( .A0(n35030), .A1(n26621), .B0(n25732), .B1(n28349), .Y(
        n25734) );
  OAI22XL U30184 ( .A0(n35033), .A1(n16672), .B0(n26246), .B1(n35239), .Y(
        n25733) );
  AOI211XL U30185 ( .A0(n16665), .A1(n26245), .B0(n25734), .C0(n25733), .Y(
        n25735) );
  NAND3XL U30186 ( .A(n25737), .B(n25736), .C(n25735), .Y(n25793) );
  OAI22XL U30187 ( .A0(n28321), .A1(n28349), .B0(n35070), .B1(n25771), .Y(
        n25742) );
  OAI22XL U30188 ( .A0(n35068), .A1(n35239), .B0(n35065), .B1(n26621), .Y(
        n25741) );
  AOI22XL U30189 ( .A0(n16665), .A1(n26199), .B0(n18463), .B1(n35069), .Y(
        n25739) );
  AOI22XL U30190 ( .A0(n35236), .A1(n35073), .B0(n16664), .B1(n26200), .Y(
        n25738) );
  OAI211XL U30191 ( .A0(n35067), .A1(n35198), .B0(n25739), .C0(n25738), .Y(
        n25740) );
  NOR3XL U30192 ( .A(n25742), .B(n25741), .C(n25740), .Y(n25780) );
  OAI22XL U30193 ( .A0(n35085), .A1(n16672), .B0(n35078), .B1(n28349), .Y(
        n25747) );
  OAI22XL U30194 ( .A0(n35081), .A1(n25771), .B0(n26223), .B1(n35200), .Y(
        n25746) );
  AOI22XL U30195 ( .A0(n35236), .A1(n35082), .B0(n16670), .B1(n26222), .Y(
        n25744) );
  AOI22XL U30196 ( .A0(n35195), .A1(n35080), .B0(n16660), .B1(n35079), .Y(
        n25743) );
  OAI211XL U30197 ( .A0(n35077), .A1(n26621), .B0(n25744), .C0(n25743), .Y(
        n25745) );
  NOR3XL U30198 ( .A(n25747), .B(n25746), .C(n25745), .Y(n25802) );
  AOI22XL U30199 ( .A0(n16670), .A1(n26192), .B0(n16664), .B1(n26191), .Y(
        n25753) );
  AOI22XL U30200 ( .A0(n35236), .A1(n35052), .B0(n25795), .B1(n35045), .Y(
        n25752) );
  OAI22XL U30201 ( .A0(n25748), .A1(n28349), .B0(n28310), .B1(n16672), .Y(
        n25750) );
  OAI22XL U30202 ( .A0(n26190), .A1(n26621), .B0(n35041), .B1(n35198), .Y(
        n25749) );
  AOI211XL U30203 ( .A0(n35195), .A1(n26193), .B0(n25750), .C0(n25749), .Y(
        n25751) );
  NAND3XL U30204 ( .A(n25753), .B(n25752), .C(n25751), .Y(n25782) );
  AOI22XL U30205 ( .A0(n35236), .A1(n35115), .B0(n18463), .B1(n25754), .Y(
        n25760) );
  AOI22XL U30206 ( .A0(n35195), .A1(n35123), .B0(n16670), .B1(n26232), .Y(
        n25759) );
  OAI22XL U30207 ( .A0(n25755), .A1(n26621), .B0(n26229), .B1(n35200), .Y(
        n25757) );
  OAI22XL U30208 ( .A0(n28339), .A1(n35198), .B0(n35112), .B1(n28349), .Y(
        n25756) );
  AOI211XL U30209 ( .A0(n25795), .A1(n35114), .B0(n25757), .C0(n25756), .Y(
        n25758) );
  NAND3XL U30210 ( .A(n25760), .B(n25759), .C(n25758), .Y(n25792) );
  OAI22XL U30211 ( .A0(n25761), .A1(n28553), .B0(n35103), .B1(n26621), .Y(
        n25765) );
  OAI22XL U30212 ( .A0(n25763), .A1(n34989), .B0(n25762), .B1(n26575), .Y(
        n25764) );
  AOI211XL U30213 ( .A0(n25766), .A1(n35104), .B0(n25765), .C0(n25764), .Y(
        n25769) );
  NAND2XL U30214 ( .A(n16664), .B(n25767), .Y(n25768) );
  OAI211XL U30215 ( .A0(n25770), .A1(n28349), .B0(n25769), .C0(n25768), .Y(
        n25779) );
  AOI22XL U30216 ( .A0(n16660), .A1(n35091), .B0(n18463), .B1(n35100), .Y(
        n25776) );
  AOI22XL U30217 ( .A0(n16670), .A1(n26215), .B0(n16664), .B1(n26214), .Y(
        n25775) );
  OAI22XL U30218 ( .A0(n35090), .A1(n25771), .B0(n26213), .B1(n18208), .Y(
        n25773) );
  OAI22XL U30219 ( .A0(n28315), .A1(n26621), .B0(n35089), .B1(n28349), .Y(
        n25772) );
  AOI211XL U30220 ( .A0(n35195), .A1(n35094), .B0(n25773), .C0(n25772), .Y(
        n25774) );
  NAND3XL U30221 ( .A(n25776), .B(n25775), .C(n25774), .Y(n25781) );
  NOR4XL U30222 ( .A(n25782), .B(n25792), .C(n25779), .D(n25781), .Y(n25777)
         );
  NAND4XL U30223 ( .A(n25778), .B(n25780), .C(n25802), .D(n25777), .Y(n25784)
         );
  INVXL U30224 ( .A(n25779), .Y(n26707) );
  OAI22XL U30225 ( .A0(n35197), .A1(n26621), .B0(n35201), .B1(n28349), .Y(
        n25790) );
  AOI22XL U30226 ( .A0(n16660), .A1(n35193), .B0(n16664), .B1(n26261), .Y(
        n25788) );
  AOI22XL U30227 ( .A0(n16670), .A1(n26259), .B0(n25795), .B1(n35206), .Y(
        n25787) );
  AOI22XL U30228 ( .A0(n35195), .A1(n28371), .B0(n18463), .B1(n28374), .Y(
        n25786) );
  NAND3XL U30229 ( .A(n25788), .B(n25787), .C(n25786), .Y(n25789) );
  AOI211XL U30230 ( .A0(n35236), .A1(n35194), .B0(n25790), .C0(n25789), .Y(
        n25791) );
  INVXL U30231 ( .A(n25791), .Y(n25803) );
  AOI22XL U30232 ( .A0(n16660), .A1(n35189), .B0(n18463), .B1(n35185), .Y(
        n25800) );
  AOI22XL U30233 ( .A0(n35195), .A1(n35180), .B0(n35236), .B1(n35179), .Y(
        n25799) );
  AOI22XL U30234 ( .A0(n16670), .A1(n26275), .B0(n25795), .B1(n28364), .Y(
        n25798) );
  OAI22XL U30235 ( .A0(n35182), .A1(n28349), .B0(n26280), .B1(n35200), .Y(
        n25796) );
  AOI2BB1XL U30236 ( .A0N(n35186), .A1N(n26621), .B0(n25796), .Y(n25797) );
  NAND4XL U30237 ( .A(n25800), .B(n25799), .C(n25798), .D(n25797), .Y(n25804)
         );
  NAND4BXL U30238 ( .AN(n25802), .B(pool[124]), .C(n25801), .D(n25804), .Y(
        n25806) );
  NOR3XL U30239 ( .A(pool[124]), .B(n25804), .C(n25803), .Y(n25805) );
  NAND2XL U30240 ( .A(n35022), .B(pool[120]), .Y(n25810) );
  OAI21XL U30241 ( .A0(n25811), .A1(n35022), .B0(n25810), .Y(N29336) );
  AOI22XL U30242 ( .A0(conv_2[239]), .A1(n26059), .B0(n25875), .B1(n25812), 
        .Y(n25830) );
  AOI22XL U30243 ( .A0(conv_2[224]), .A1(n26082), .B0(n26081), .B1(n25813), 
        .Y(n25829) );
  OAI22XL U30244 ( .A0(n35143), .A1(n25816), .B0(n28479), .B1(n25815), .Y(
        n25817) );
  AOI211XL U30245 ( .A0(n34903), .A1(n25819), .B0(n25818), .C0(n25817), .Y(
        n25828) );
  OAI22XL U30246 ( .A0(n25821), .A1(n18208), .B0(n25820), .B1(n26039), .Y(
        n25825) );
  OAI22XL U30247 ( .A0(n25823), .A1(n35198), .B0(n25822), .B1(n35239), .Y(
        n25824) );
  AOI211XL U30248 ( .A0(n16755), .A1(n25826), .B0(n25825), .C0(n25824), .Y(
        n25827) );
  NAND4XL U30249 ( .A(n25830), .B(n25829), .C(n25828), .D(n25827), .Y(n26111)
         );
  OAI2BB1XL U30250 ( .A0N(n35231), .A1N(n25831), .B0(n26026), .Y(n25832) );
  AOI22XL U30251 ( .A0(n35236), .A1(n25834), .B0(n25833), .B1(n25832), .Y(
        n25835) );
  OAI21XL U30252 ( .A0(n25836), .A1(n25987), .B0(n25835), .Y(n25848) );
  AOI22XL U30253 ( .A0(conv_2[228]), .A1(n26059), .B0(n34903), .B1(n25837), 
        .Y(n25846) );
  AOI22XL U30254 ( .A0(n26082), .A1(conv_2[213]), .B0(n26081), .B1(n25838), 
        .Y(n25845) );
  AOI22XL U30255 ( .A0(n16660), .A1(n25840), .B0(n19179), .B1(n25839), .Y(
        n25844) );
  AOI22XL U30256 ( .A0(n35195), .A1(n25842), .B0(n16671), .B1(n25841), .Y(
        n25843) );
  NAND4XL U30257 ( .A(n25846), .B(n25845), .C(n25844), .D(n25843), .Y(n25847)
         );
  AOI22XL U30258 ( .A0(conv_2[212]), .A1(n26082), .B0(n16671), .B1(n25850), 
        .Y(n25851) );
  OAI21XL U30259 ( .A0(n25853), .A1(n25852), .B0(n25851), .Y(n25866) );
  AOI22XL U30260 ( .A0(conv_2[227]), .A1(n26059), .B0(n26066), .B1(n25854), 
        .Y(n25864) );
  AOI22XL U30261 ( .A0(n19179), .A1(n25856), .B0(n34903), .B1(n25855), .Y(
        n25863) );
  AOI22XL U30262 ( .A0(n35195), .A1(n25858), .B0(n34906), .B1(n25857), .Y(
        n25862) );
  AOI22XL U30263 ( .A0(n35236), .A1(n25860), .B0(n16660), .B1(n25859), .Y(
        n25861) );
  NAND4XL U30264 ( .A(n25864), .B(n25863), .C(n25862), .D(n25861), .Y(n25865)
         );
  AOI22XL U30265 ( .A0(n16660), .A1(n25870), .B0(conv_2[211]), .B1(n26082), 
        .Y(n25871) );
  OAI21XL U30266 ( .A0(n25873), .A1(n25872), .B0(n25871), .Y(n25888) );
  AOI22XL U30267 ( .A0(n34903), .A1(n25876), .B0(n25875), .B1(n25874), .Y(
        n25886) );
  AOI22XL U30268 ( .A0(n35195), .A1(n25877), .B0(conv_2[226]), .B1(n26059), 
        .Y(n25885) );
  AOI22XL U30269 ( .A0(n35236), .A1(n25880), .B0(n25879), .B1(n25878), .Y(
        n25884) );
  AOI22XL U30270 ( .A0(n19179), .A1(n25882), .B0(n16671), .B1(n25881), .Y(
        n25883) );
  NAND4XL U30271 ( .A(n25886), .B(n25885), .C(n25884), .D(n25883), .Y(n25887)
         );
  AOI222XL U30272 ( .A0(pool[80]), .A1(pool[81]), .B0(pool[80]), .B1(n26113), 
        .C0(pool[81]), .C1(n26113), .Y(n25890) );
  AOI222XL U30273 ( .A0(n34925), .A1(n34924), .B0(n34925), .B1(n25890), .C0(
        n34924), .C1(n25890), .Y(n25891) );
  AOI222XL U30274 ( .A0(n26118), .A1(pool[83]), .B0(n26118), .B1(n25891), .C0(
        pool[83]), .C1(n25891), .Y(n26057) );
  AOI22XL U30275 ( .A0(conv_2[230]), .A1(n26059), .B0(n26276), .B1(n25892), 
        .Y(n25895) );
  NAND2XL U30276 ( .A(n16671), .B(n25893), .Y(n25894) );
  OAI211XL U30277 ( .A0(n35143), .A1(n25896), .B0(n25895), .C0(n25894), .Y(
        n25909) );
  AOI22XL U30278 ( .A0(n26082), .A1(conv_2[215]), .B0(n34903), .B1(n25897), 
        .Y(n25907) );
  AOI22XL U30279 ( .A0(n28528), .A1(n25899), .B0(n26081), .B1(n25898), .Y(
        n25906) );
  AOI22XL U30280 ( .A0(n16660), .A1(n25901), .B0(n19179), .B1(n25900), .Y(
        n25905) );
  AOI22XL U30281 ( .A0(n35195), .A1(n25903), .B0(n35236), .B1(n25902), .Y(
        n25904) );
  NAND4XL U30282 ( .A(n25907), .B(n25906), .C(n25905), .D(n25904), .Y(n25908)
         );
  AOI211XL U30283 ( .A0(n16755), .A1(n25910), .B0(n25909), .C0(n25908), .Y(
        n26053) );
  AOI22XL U30284 ( .A0(n26059), .A1(conv_2[232]), .B0(n26081), .B1(n25911), 
        .Y(n25914) );
  NAND2XL U30285 ( .A(n26066), .B(n25912), .Y(n25913) );
  OAI211XL U30286 ( .A0(n25915), .A1(n26026), .B0(n25914), .C0(n25913), .Y(
        n25928) );
  AOI22XL U30287 ( .A0(n16660), .A1(n25916), .B0(conv_2[217]), .B1(n26082), 
        .Y(n25926) );
  AOI22XL U30288 ( .A0(n34903), .A1(n25918), .B0(n35231), .B1(n25917), .Y(
        n25925) );
  AOI22XL U30289 ( .A0(n35195), .A1(n25920), .B0(n35236), .B1(n25919), .Y(
        n25924) );
  AOI22XL U30290 ( .A0(n19179), .A1(n25922), .B0(n16671), .B1(n25921), .Y(
        n25923) );
  NAND4XL U30291 ( .A(n25926), .B(n25925), .C(n25924), .D(n25923), .Y(n25927)
         );
  AOI211XL U30292 ( .A0(n16755), .A1(n25929), .B0(n25928), .C0(n25927), .Y(
        n26052) );
  INVXL U30293 ( .A(conv_2[229]), .Y(n29054) );
  AOI22XL U30294 ( .A0(n35236), .A1(n25931), .B0(n26081), .B1(n25930), .Y(
        n25948) );
  AOI22XL U30295 ( .A0(conv_2[214]), .A1(n26082), .B0(n16671), .B1(n25932), 
        .Y(n25935) );
  NAND2XL U30296 ( .A(n16660), .B(n25933), .Y(n25934) );
  OAI211XL U30297 ( .A0(n25936), .A1(n26026), .B0(n25935), .C0(n25934), .Y(
        n25945) );
  AOI22XL U30298 ( .A0(n35195), .A1(n25938), .B0(n19179), .B1(n25937), .Y(
        n25942) );
  OAI21XL U30299 ( .A0(n25940), .A1(n25939), .B0(n28528), .Y(n25941) );
  OAI211XL U30300 ( .A0(n35143), .A1(n25943), .B0(n25942), .C0(n25941), .Y(
        n25944) );
  AOI211XL U30301 ( .A0(n16755), .A1(n25946), .B0(n25945), .C0(n25944), .Y(
        n25947) );
  OAI211XL U30302 ( .A0(n29054), .A1(n26085), .B0(n25948), .C0(n25947), .Y(
        n26051) );
  AOI22XL U30303 ( .A0(n16671), .A1(n25950), .B0(n26081), .B1(n25949), .Y(
        n25968) );
  AOI22XL U30304 ( .A0(n35236), .A1(n25952), .B0(n18197), .B1(n25951), .Y(
        n25954) );
  NAND2XL U30305 ( .A(conv_2[216]), .B(n26082), .Y(n25953) );
  OAI211XL U30306 ( .A0(n25955), .A1(n26026), .B0(n25954), .C0(n25953), .Y(
        n25965) );
  AOI22XL U30307 ( .A0(n19179), .A1(n25957), .B0(n25956), .B1(n35231), .Y(
        n25962) );
  OAI211XL U30308 ( .A0(n25963), .A1(n35239), .B0(n25962), .C0(n25961), .Y(
        n25964) );
  AOI211XL U30309 ( .A0(n16755), .A1(n25966), .B0(n25965), .C0(n25964), .Y(
        n25967) );
  OAI211XL U30310 ( .A0(n29178), .A1(n26085), .B0(n25968), .C0(n25967), .Y(
        n26054) );
  AOI22XL U30311 ( .A0(n16660), .A1(n25970), .B0(n26081), .B1(n25969), .Y(
        n25986) );
  AOI22XL U30312 ( .A0(n19179), .A1(n25972), .B0(n16671), .B1(n25971), .Y(
        n25973) );
  OAI21XL U30313 ( .A0(n25975), .A1(n25974), .B0(n25973), .Y(n25983) );
  AOI22XL U30314 ( .A0(conv_2[218]), .A1(n26082), .B0(n34903), .B1(n25976), 
        .Y(n25980) );
  AOI22XL U30315 ( .A0(n35195), .A1(n25978), .B0(n26276), .B1(n25977), .Y(
        n25979) );
  OAI211XL U30316 ( .A0(n25981), .A1(n35159), .B0(n25980), .C0(n25979), .Y(
        n25982) );
  AOI211XL U30317 ( .A0(n35236), .A1(n25984), .B0(n25983), .C0(n25982), .Y(
        n25985) );
  OAI211XL U30318 ( .A0(n29188), .A1(n26085), .B0(n25986), .C0(n25985), .Y(
        n26101) );
  OAI22XL U30319 ( .A0(n30429), .A1(n26029), .B0(n35196), .B1(n25989), .Y(
        n25990) );
  AOI211XL U30320 ( .A0(n34903), .A1(n25992), .B0(n25991), .C0(n25990), .Y(
        n26006) );
  AOI22XL U30321 ( .A0(n19179), .A1(n25994), .B0(n35231), .B1(n25993), .Y(
        n26005) );
  AOI22XL U30322 ( .A0(n35195), .A1(n25996), .B0(n16671), .B1(n25995), .Y(
        n26004) );
  OAI22XL U30323 ( .A0(n25997), .A1(n26026), .B0(n29159), .B1(n26085), .Y(
        n26001) );
  OAI22XL U30324 ( .A0(n25999), .A1(n35198), .B0(n25998), .B1(n18208), .Y(
        n26000) );
  AOI211XL U30325 ( .A0(n16755), .A1(n26002), .B0(n26001), .C0(n26000), .Y(
        n26003) );
  NAND4XL U30326 ( .A(n26006), .B(n26005), .C(n26004), .D(n26003), .Y(n26104)
         );
  AOI22XL U30327 ( .A0(n16660), .A1(n26008), .B0(n26081), .B1(n26007), .Y(
        n26025) );
  AOI22XL U30328 ( .A0(conv_2[221]), .A1(n26082), .B0(conv_2[236]), .B1(n26059), .Y(n26013) );
  OAI211XL U30329 ( .A0(n26014), .A1(n18208), .B0(n26013), .C0(n26012), .Y(
        n26023) );
  AOI22XL U30330 ( .A0(n19179), .A1(n26016), .B0(n26015), .B1(n35231), .Y(
        n26020) );
  AOI22XL U30331 ( .A0(n35195), .A1(n26018), .B0(n16671), .B1(n26017), .Y(
        n26019) );
  OAI211XL U30332 ( .A0(n26021), .A1(n35159), .B0(n26020), .C0(n26019), .Y(
        n26022) );
  OAI211XL U30333 ( .A0(n26027), .A1(n26026), .B0(n26025), .C0(n26024), .Y(
        n26103) );
  OAI22XL U30334 ( .A0(n30434), .A1(n26029), .B0(n26162), .B1(n26028), .Y(
        n26030) );
  AOI211XL U30335 ( .A0(n26081), .A1(n26032), .B0(n26031), .C0(n26030), .Y(
        n26048) );
  AOI22XL U30336 ( .A0(n16660), .A1(n26034), .B0(n35231), .B1(n26033), .Y(
        n26047) );
  AOI22XL U30337 ( .A0(n35236), .A1(n26036), .B0(n16671), .B1(n26035), .Y(
        n26046) );
  OAI22XL U30338 ( .A0(n26038), .A1(n26086), .B0(n28479), .B1(n26037), .Y(
        n26043) );
  OAI22XL U30339 ( .A0(n26041), .A1(n35239), .B0(n26040), .B1(n26039), .Y(
        n26042) );
  AOI211XL U30340 ( .A0(n16755), .A1(n26044), .B0(n26043), .C0(n26042), .Y(
        n26045) );
  NAND4XL U30341 ( .A(n26048), .B(n26047), .C(n26046), .D(n26045), .Y(n26102)
         );
  NOR4XL U30342 ( .A(n26101), .B(n26104), .C(n26103), .D(n26102), .Y(n26049)
         );
  NAND4XL U30343 ( .A(n26053), .B(n26052), .C(n26050), .D(n26049), .Y(n26056)
         );
  INVXL U30344 ( .A(n26051), .Y(n26115) );
  AOI22XL U30345 ( .A0(conv_2[237]), .A1(n26059), .B0(n16671), .B1(n26058), 
        .Y(n26062) );
  NAND2XL U30346 ( .A(n19179), .B(n26060), .Y(n26061) );
  OAI211XL U30347 ( .A0(n26162), .A1(n26063), .B0(n26062), .C0(n26061), .Y(
        n26077) );
  AOI22XL U30348 ( .A0(n26066), .A1(n26065), .B0(n26081), .B1(n26064), .Y(
        n26075) );
  AOI22XL U30349 ( .A0(conv_2[222]), .A1(n26082), .B0(n34903), .B1(n26067), 
        .Y(n26074) );
  AOI22XL U30350 ( .A0(n35195), .A1(n26069), .B0(n35236), .B1(n26068), .Y(
        n26073) );
  AOI22XL U30351 ( .A0(n16660), .A1(n26071), .B0(n35231), .B1(n26070), .Y(
        n26072) );
  NAND4XL U30352 ( .A(n26075), .B(n26074), .C(n26073), .D(n26072), .Y(n26076)
         );
  AOI211XL U30353 ( .A0(n16755), .A1(n26078), .B0(n26077), .C0(n26076), .Y(
        n26079) );
  INVXL U30354 ( .A(n26079), .Y(n26106) );
  AOI22XL U30355 ( .A0(conv_2[223]), .A1(n26082), .B0(n26081), .B1(n26080), 
        .Y(n26084) );
  AOI32XL U30356 ( .A0(n35143), .A1(n26084), .A2(n26162), .B0(n26083), .B1(
        n26084), .Y(n26100) );
  OAI22XL U30357 ( .A0(n26087), .A1(n26086), .B0(n26085), .B1(n33094), .Y(
        n26099) );
  OAI22XL U30358 ( .A0(n35184), .A1(n26089), .B0(n26088), .B1(n18208), .Y(
        n26098) );
  AOI22XL U30359 ( .A0(n16660), .A1(n26091), .B0(n16671), .B1(n26090), .Y(
        n26095) );
  AOI22XL U30360 ( .A0(n35195), .A1(n26093), .B0(n19179), .B1(n26092), .Y(
        n26094) );
  OAI211XL U30361 ( .A0(n26096), .A1(n35159), .B0(n26095), .C0(n26094), .Y(
        n26097) );
  NAND4XL U30362 ( .A(n26105), .B(n26104), .C(n26103), .D(n26102), .Y(n26109)
         );
  NOR3XL U30363 ( .A(pool[84]), .B(n26107), .C(n26106), .Y(n26108) );
  INVXL U30364 ( .A(n34926), .Y(n26117) );
  AOI22XL U30365 ( .A0(n34926), .A1(n26114), .B0(n26113), .B1(n26117), .Y(
        N29297) );
  AOI22XL U30366 ( .A0(n34926), .A1(n26116), .B0(n26115), .B1(n26117), .Y(
        N29300) );
  AOI22XL U30367 ( .A0(n34926), .A1(n26119), .B0(n26118), .B1(n26117), .Y(
        N29299) );
  OAI21XL U30368 ( .A0(n26123), .A1(n16654), .B0(n35813), .Y(n26122) );
  NAND2XL U30369 ( .A(n26125), .B(n35588), .Y(n15433) );
  INVXL U30370 ( .A(conv_1[56]), .Y(n29753) );
  NAND2XL U30371 ( .A(n27230), .B(n34507), .Y(n26131) );
  INVXL U30372 ( .A(conv_1[45]), .Y(n33514) );
  AOI2BB1XL U30373 ( .A0N(n35272), .A1N(n27799), .B0(n33512), .Y(n26126) );
  INVXL U30374 ( .A(n26126), .Y(n27467) );
  NAND2XL U30375 ( .A(n33512), .B(n27429), .Y(n27466) );
  NAND2XL U30376 ( .A(n27471), .B(n27466), .Y(n26127) );
  NAND2XL U30377 ( .A(n27467), .B(n26127), .Y(n26128) );
  OAI21XL U30378 ( .A0(n33403), .A1(n27799), .B0(n26128), .Y(n26129) );
  INVXL U30379 ( .A(n26129), .Y(n27439) );
  AOI222XL U30380 ( .A0(n27327), .A1(n27326), .B0(n27327), .B1(conv_1[48]), 
        .C0(n27326), .C1(conv_1[48]), .Y(n26130) );
  NOR2X1 U30381 ( .A(n26131), .B(n26130), .Y(n27456) );
  NAND2XL U30382 ( .A(n35316), .B(n26133), .Y(n26132) );
  OAI21XL U30383 ( .A0(conv_1[55]), .A1(n35314), .B0(n35316), .Y(n29752) );
  INVXL U30384 ( .A(conv_1[52]), .Y(n26824) );
  NAND2XL U30385 ( .A(conv_1[50]), .B(n27323), .Y(n27322) );
  NAND2XL U30386 ( .A(conv_1[51]), .B(n27313), .Y(n27312) );
  NAND2XL U30387 ( .A(conv_1[53]), .B(n27317), .Y(n35308) );
  OAI2BB1XL U30388 ( .A0N(conv_1[55]), .A1N(n35315), .B0(n35309), .Y(n32517)
         );
  NAND2XL U30389 ( .A(n29752), .B(n32517), .Y(n26136) );
  AOI211XL U30390 ( .A0(n29753), .A1(n26136), .B0(n36042), .C0(n26135), .Y(
        n26137) );
  AOI2BB1XL U30391 ( .A0N(n29753), .A1N(n35319), .B0(n26137), .Y(n26138) );
  NAND2XL U30392 ( .A(n26138), .B(n34544), .Y(n16407) );
  INVXL U30393 ( .A(n35324), .Y(n33638) );
  ADDFX1 U30394 ( .A(conv_1[63]), .B(n26140), .CI(n26139), .CO(n27406), .S(
        n22420) );
  AOI222XL U30395 ( .A0(n27405), .A1(n27406), .B0(n27405), .B1(conv_1[64]), 
        .C0(n27406), .C1(conv_1[64]), .Y(n26141) );
  INVXL U30396 ( .A(conv_1[67]), .Y(n35326) );
  INVXL U30397 ( .A(conv_1[65]), .Y(n27111) );
  NAND2XL U30398 ( .A(conv_1[66]), .B(n27101), .Y(n35323) );
  NAND2XL U30399 ( .A(conv_1[68]), .B(n27201), .Y(n27095) );
  AOI21XL U30400 ( .A0(conv_1[70]), .A1(n33637), .B0(n33638), .Y(n27088) );
  AOI22XL U30401 ( .A0(n33638), .A1(n26311), .B0(n26309), .B1(n35324), .Y(
        n26143) );
  AOI211XL U30402 ( .A0(n26310), .A1(n26143), .B0(n36009), .C0(n26142), .Y(
        n26144) );
  NAND2XL U30403 ( .A(n26145), .B(n34281), .Y(n16391) );
  OAI21XL U30404 ( .A0(n16654), .A1(n26146), .B0(n33432), .Y(n26147) );
  AOI22XL U30405 ( .A0(n32660), .A1(n26148), .B0(conv_1[529]), .B1(n26147), 
        .Y(n26149) );
  NAND2XL U30406 ( .A(n26149), .B(n35489), .Y(n15934) );
  AOI22XL U30407 ( .A0(n34884), .A1(n26151), .B0(n26150), .B1(n34885), .Y(
        N29280) );
  OAI21XL U30408 ( .A0(n26156), .A1(n16655), .B0(n35676), .Y(n26155) );
  AOI32XL U30409 ( .A0(n36020), .A1(n29160), .A2(n26156), .B0(conv_3[230]), 
        .B1(n26155), .Y(n26157) );
  NAND2XL U30410 ( .A(n26157), .B(n35588), .Y(n15593) );
  OAI22XL U30411 ( .A0(n34982), .A1(n26207), .B0(n35240), .B1(n28479), .Y(
        n26161) );
  AOI22XL U30412 ( .A0(n26263), .A1(n35232), .B0(n16667), .B1(n35235), .Y(
        n26158) );
  OAI21XL U30413 ( .A0(n26159), .A1(n28467), .B0(n26158), .Y(n26160) );
  AOI22XL U30414 ( .A0(n26263), .A1(n35167), .B0(n16667), .B1(n28264), .Y(
        n26169) );
  OAI22XL U30415 ( .A0(n26163), .A1(n26162), .B0(n35171), .B1(n26274), .Y(
        n26165) );
  OAI2BB2XL U30416 ( .B0(n35170), .B1(n26285), .A0N(n35168), .A1N(n28528), .Y(
        n26164) );
  AOI211XL U30417 ( .A0(n26262), .A1(n26166), .B0(n26165), .C0(n26164), .Y(
        n26167) );
  NAND3XL U30418 ( .A(n26169), .B(n26168), .C(n26167), .Y(n26293) );
  AOI22XL U30419 ( .A0(n16667), .A1(n35127), .B0(n26172), .B1(n26171), .Y(
        n26173) );
  OAI211XL U30420 ( .A0(n26175), .A1(n28467), .B0(n26174), .C0(n26173), .Y(
        n26176) );
  AOI21XL U30421 ( .A0(n28467), .A1(n16721), .B0(n26177), .Y(n26181) );
  AOI22XL U30422 ( .A0(n26263), .A1(n35151), .B0(n16667), .B1(n35154), .Y(
        n26178) );
  AOI211XL U30423 ( .A0(n28528), .A1(n35152), .B0(n26181), .C0(n26180), .Y(
        n27069) );
  AOI222XL U30424 ( .A0(pool[91]), .A1(n26296), .B0(pool[91]), .B1(n27069), 
        .C0(n26296), .C1(n27069), .Y(n26188) );
  AOI22XL U30425 ( .A0(n26263), .A1(n26182), .B0(n16667), .B1(n35140), .Y(
        n26187) );
  NAND2XL U30426 ( .A(n36244), .B(n28278), .Y(n26185) );
  NAND2XL U30427 ( .A(n28528), .B(n35148), .Y(n26184) );
  NAND4XL U30428 ( .A(n26187), .B(n26186), .C(n26185), .D(n26184), .Y(n34944)
         );
  INVXL U30429 ( .A(pool[92]), .Y(n34946) );
  AOI222XL U30430 ( .A0(n26188), .A1(n34944), .B0(n26188), .B1(n34946), .C0(
        n34944), .C1(n34946), .Y(n26189) );
  AOI222XL U30431 ( .A0(pool[93]), .A1(n34947), .B0(pool[93]), .B1(n26189), 
        .C0(n34947), .C1(n26189), .Y(n26258) );
  INVXL U30432 ( .A(pool[94]), .Y(n27066) );
  OAI22XL U30433 ( .A0(n28310), .A1(n16661), .B0(n35041), .B1(n28577), .Y(
        n26198) );
  INVXL U30434 ( .A(n26190), .Y(n35044) );
  AOI22XL U30435 ( .A0(n26262), .A1(n26191), .B0(n26260), .B1(n35044), .Y(
        n26196) );
  AOI22XL U30436 ( .A0(n26376), .A1(n35043), .B0(n26276), .B1(n26192), .Y(
        n26195) );
  NAND3XL U30437 ( .A(n26196), .B(n26195), .C(n26194), .Y(n26197) );
  AOI211XL U30438 ( .A0(n36244), .A1(n35045), .B0(n26198), .C0(n26197), .Y(
        n26252) );
  OAI22XL U30439 ( .A0(n28321), .A1(n26274), .B0(n35070), .B1(n16721), .Y(
        n26205) );
  OAI22XL U30440 ( .A0(n35065), .A1(n26285), .B0(n35067), .B1(n28577), .Y(
        n26204) );
  AOI22XL U30441 ( .A0(n26262), .A1(n26200), .B0(n26276), .B1(n26199), .Y(
        n26202) );
  AOI22XL U30442 ( .A0(n26263), .A1(n35069), .B0(n28528), .B1(n35073), .Y(
        n26201) );
  NAND2XL U30443 ( .A(n26202), .B(n26201), .Y(n26203) );
  NOR4XL U30444 ( .A(n26206), .B(n26205), .C(n26204), .D(n26203), .Y(n26253)
         );
  OAI22XL U30445 ( .A0(n24828), .A1(n26207), .B0(n35107), .B1(n28479), .Y(
        n26212) );
  OAI21XL U30446 ( .A0(n26210), .A1(n28467), .B0(n26209), .Y(n26211) );
  OAI22XL U30447 ( .A0(n35090), .A1(n16721), .B0(n26213), .B1(n28479), .Y(
        n26221) );
  AOI22XL U30448 ( .A0(n16667), .A1(n35091), .B0(n26262), .B1(n26214), .Y(
        n26219) );
  AOI22XL U30449 ( .A0(n26260), .A1(n35093), .B0(n26276), .B1(n26215), .Y(
        n26218) );
  AOI22XL U30450 ( .A0(n26263), .A1(n35100), .B0(n26376), .B1(n26216), .Y(
        n26217) );
  NAND3XL U30451 ( .A(n26219), .B(n26218), .C(n26217), .Y(n26220) );
  AOI22XL U30452 ( .A0(n16667), .A1(n35079), .B0(n26276), .B1(n26222), .Y(
        n26228) );
  INVXL U30453 ( .A(n35080), .Y(n28331) );
  OAI22XL U30454 ( .A0(n35078), .A1(n26274), .B0(n28331), .B1(n28575), .Y(
        n26226) );
  OAI22XL U30455 ( .A0(n26223), .A1(n26279), .B0(n35077), .B1(n26285), .Y(
        n26225) );
  OAI22XL U30456 ( .A0(n35085), .A1(n34958), .B0(n28332), .B1(n28479), .Y(
        n26224) );
  NOR3XL U30457 ( .A(n26226), .B(n26225), .C(n26224), .Y(n26227) );
  OAI211XL U30458 ( .A0(n35081), .A1(n16721), .B0(n26228), .C0(n26227), .Y(
        n26272) );
  AOI22XL U30459 ( .A0(n36244), .A1(n35114), .B0(n26260), .B1(n35116), .Y(
        n26235) );
  OAI22XL U30460 ( .A0(n35113), .A1(n34958), .B0(n28339), .B1(n28577), .Y(
        n26231) );
  OAI22XL U30461 ( .A0(n26229), .A1(n26279), .B0(n35112), .B1(n26274), .Y(
        n26230) );
  AOI211XL U30462 ( .A0(n26276), .A1(n26232), .B0(n26231), .C0(n26230), .Y(
        n26233) );
  NAND3XL U30463 ( .A(n26235), .B(n26234), .C(n26233), .Y(n26271) );
  AOI22XL U30464 ( .A0(n36244), .A1(n35054), .B0(n26376), .B1(n28352), .Y(
        n26243) );
  AOI22XL U30465 ( .A0(n28528), .A1(n35061), .B0(n26262), .B1(n26237), .Y(
        n26242) );
  OAI22XL U30466 ( .A0(n35058), .A1(n28577), .B0(n35055), .B1(n28575), .Y(
        n26239) );
  OAI22XL U30467 ( .A0(n35053), .A1(n26285), .B0(n35057), .B1(n34958), .Y(
        n26238) );
  AOI211XL U30468 ( .A0(n26276), .A1(n26240), .B0(n26239), .C0(n26238), .Y(
        n26241) );
  NAND3XL U30469 ( .A(n26243), .B(n26242), .C(n26241), .Y(n26286) );
  AOI22XL U30470 ( .A0(n26376), .A1(n35031), .B0(n26262), .B1(n26244), .Y(
        n26251) );
  AOI22XL U30471 ( .A0(n36244), .A1(n35034), .B0(n26276), .B1(n26245), .Y(
        n26250) );
  OAI22XL U30472 ( .A0(n35033), .A1(n34958), .B0(n26246), .B1(n28575), .Y(
        n26248) );
  INVXL U30473 ( .A(n28344), .Y(n35029) );
  OAI22XL U30474 ( .A0(n35030), .A1(n26285), .B0(n35029), .B1(n28577), .Y(
        n26247) );
  AOI211XL U30475 ( .A0(n28528), .A1(n35040), .B0(n26248), .C0(n26247), .Y(
        n26249) );
  NAND3XL U30476 ( .A(n26251), .B(n26250), .C(n26249), .Y(n26273) );
  NOR4BBXL U30477 ( .AN(n26253), .BN(n26252), .C(n26286), .D(n26273), .Y(
        n26254) );
  NAND2XL U30478 ( .A(n26255), .B(n26254), .Y(n26256) );
  AOI22XL U30479 ( .A0(n26260), .A1(n28373), .B0(n26276), .B1(n26259), .Y(
        n26267) );
  AOI22XL U30480 ( .A0(n26263), .A1(n28374), .B0(n28528), .B1(n35194), .Y(
        n26265) );
  NAND2XL U30481 ( .A(n28556), .B(n35193), .Y(n26264) );
  NAND4XL U30482 ( .A(n26267), .B(n26266), .C(n26265), .D(n26264), .Y(n26268)
         );
  AOI211XL U30483 ( .A0(n36244), .A1(n35206), .B0(n26269), .C0(n26268), .Y(
        n26270) );
  INVXL U30484 ( .A(n26270), .Y(n26288) );
  AOI22XL U30485 ( .A0(n28556), .A1(n35189), .B0(n26276), .B1(n26275), .Y(
        n26278) );
  AOI22XL U30486 ( .A0(n36244), .A1(n28364), .B0(n26263), .B1(n35185), .Y(
        n26277) );
  OAI211XL U30487 ( .A0(n26280), .A1(n26279), .B0(n26278), .C0(n26277), .Y(
        n26281) );
  NAND2XL U30488 ( .A(n28528), .B(n35179), .Y(n26283) );
  OAI211XL U30489 ( .A0(n35186), .A1(n26285), .B0(n26284), .C0(n26283), .Y(
        n26289) );
  NAND4XL U30490 ( .A(pool[94]), .B(n26287), .C(n26289), .D(n26286), .Y(n26291) );
  NOR3XL U30491 ( .A(pool[94]), .B(n26289), .C(n26288), .Y(n26290) );
  NAND2XL U30492 ( .A(n34945), .B(pool[90]), .Y(n26295) );
  OAI21XL U30493 ( .A0(n26296), .A1(n34945), .B0(n26295), .Y(N29306) );
  NAND2XL U30494 ( .A(n26297), .B(n34547), .Y(n27364) );
  NAND2XL U30495 ( .A(n27364), .B(n27363), .Y(n26300) );
  OAI21XL U30496 ( .A0(n16654), .A1(n26300), .B0(n34552), .Y(n26299) );
  NAND2XL U30497 ( .A(n26301), .B(n34682), .Y(n16450) );
  ADDFXL U30498 ( .A(conv_3[530]), .B(n33719), .CI(n26302), .CO(n26369), .S(
        n24366) );
  NAND2XL U30499 ( .A(n33719), .B(n26369), .Y(n26303) );
  OAI21XL U30500 ( .A0(n33719), .A1(n26369), .B0(n26303), .Y(n26305) );
  AOI211XL U30501 ( .A0(n26307), .A1(n26305), .B0(n16658), .C0(n26304), .Y(
        n26306) );
  AOI2BB1XL U30502 ( .A0N(n26307), .A1N(n31191), .B0(n26306), .Y(n26308) );
  NAND2XL U30503 ( .A(n26308), .B(n35588), .Y(n15392) );
  INVXL U30504 ( .A(conv_1[73]), .Y(n27205) );
  NAND3XL U30505 ( .A(n26309), .B(conv_1[72]), .C(n35324), .Y(n27207) );
  NAND3XL U30506 ( .A(n26311), .B(n33638), .C(n26310), .Y(n27206) );
  NAND2XL U30507 ( .A(n27207), .B(n27206), .Y(n26313) );
  OAI21XL U30508 ( .A0(n16654), .A1(n26313), .B0(n35327), .Y(n26312) );
  AOI32XL U30509 ( .A0(n16657), .A1(n27205), .A2(n26313), .B0(conv_1[73]), 
        .B1(n26312), .Y(n26314) );
  NAND2XL U30510 ( .A(n26314), .B(n34281), .Y(n16390) );
  INVXL U30511 ( .A(n32649), .Y(n32207) );
  NOR2X1 U30512 ( .A(n32649), .B(n26317), .Y(n31615) );
  INVXL U30513 ( .A(conv_3[187]), .Y(n31601) );
  NAND2XL U30514 ( .A(n32207), .B(n31609), .Y(n26318) );
  INVXL U30515 ( .A(n26318), .Y(n26322) );
  OAI31XL U30516 ( .A0(conv_3[187]), .A1(n31597), .A2(conv_3[188]), .B0(n32649), .Y(n26319) );
  NAND2X1 U30517 ( .A(n31608), .B(n26319), .Y(n31607) );
  AOI32XL U30518 ( .A0(n26319), .A1(n34704), .A2(n26318), .B0(n34389), .B1(
        n34704), .Y(n26320) );
  AOI21XL U30519 ( .A0(conv_3[189]), .A1(n26320), .B0(n16653), .Y(n26321) );
  OAI31XL U30520 ( .A0(n26322), .A1(n16655), .A2(n31607), .B0(n26321), .Y(
        n15619) );
  INVXL U30521 ( .A(conv_1[430]), .Y(n26325) );
  INVXL U30522 ( .A(conv_1[428]), .Y(n27585) );
  NAND2XL U30523 ( .A(conv_1[427]), .B(n29402), .Y(n27584) );
  AOI21XL U30524 ( .A0(conv_1[429]), .A1(n33394), .B0(intadd_1_B_2_), .Y(
        n29222) );
  OAI21XL U30525 ( .A0(n26324), .A1(n16654), .B0(n35504), .Y(n26323) );
  AOI32XL U30526 ( .A0(n32660), .A1(n26325), .A2(n26324), .B0(conv_1[430]), 
        .B1(n26323), .Y(n26326) );
  NAND2XL U30527 ( .A(n26326), .B(n34689), .Y(n16033) );
  OAI21XL U30528 ( .A0(conv_3[274]), .A1(n26328), .B0(n26327), .Y(n26329) );
  NAND2XL U30529 ( .A(n32599), .B(n26329), .Y(n31733) );
  OR2XL U30530 ( .A(n32599), .B(n26329), .Y(n31731) );
  NAND2XL U30531 ( .A(n31733), .B(n31731), .Y(n26331) );
  AOI211XL U30532 ( .A0(n31732), .A1(n26331), .B0(n36001), .C0(n26330), .Y(
        n26332) );
  AOI2BB1XL U30533 ( .A0N(n31732), .A1N(n34709), .B0(n26332), .Y(n26333) );
  NAND2XL U30534 ( .A(n26333), .B(n35588), .Y(n15563) );
  OAI21XL U30535 ( .A0(n27131), .A1(n26335), .B0(n26334), .Y(n26337) );
  AOI211XL U30536 ( .A0(n26339), .A1(n26337), .B0(n16655), .C0(n26336), .Y(
        n26338) );
  AOI2BB1XL U30537 ( .A0N(n26339), .A1N(n33427), .B0(n26338), .Y(n26340) );
  NAND2XL U30538 ( .A(n26340), .B(n34682), .Y(n15962) );
  NAND2BXL U30539 ( .AN(n26342), .B(n26341), .Y(n26344) );
  AOI211XL U30540 ( .A0(n26346), .A1(n26344), .B0(n16655), .C0(n26343), .Y(
        n26345) );
  AOI2BB1XL U30541 ( .A0N(n26346), .A1N(n33506), .B0(n26345), .Y(n26347) );
  NAND2XL U30542 ( .A(n26347), .B(n34281), .Y(n15989) );
  AOI22XL U30543 ( .A0(n34896), .A1(n26349), .B0(n26348), .B1(n34892), .Y(
        N29290) );
  AOI22XL U30544 ( .A0(n34896), .A1(n26351), .B0(n26350), .B1(n34892), .Y(
        N29289) );
  INVXL U30545 ( .A(n35982), .Y(n33079) );
  INVXL U30546 ( .A(conv_2[322]), .Y(n35985) );
  NAND2XL U30547 ( .A(conv_2[323]), .B(n28045), .Y(n28056) );
  OAI31XL U30548 ( .A0(conv_2[322]), .A1(conv_2[323]), .A2(n35983), .B0(n35982), .Y(n28057) );
  OAI2BB1XL U30549 ( .A0N(n33079), .A1N(n28056), .B0(n28057), .Y(n26354) );
  AOI211XL U30550 ( .A0(n28058), .A1(n26354), .B0(n16655), .C0(n26353), .Y(
        n26355) );
  AOI2BB1XL U30551 ( .A0N(n28058), .A1N(n35986), .B0(n26355), .Y(n26356) );
  NAND2XL U30552 ( .A(n26356), .B(n35859), .Y(n14989) );
  OAI21XL U30553 ( .A0(n16654), .A1(n26360), .B0(n34631), .Y(n26359) );
  NAND2XL U30554 ( .A(n26362), .B(n35859), .Y(n15095) );
  OAI21XL U30555 ( .A0(n26366), .A1(n16654), .B0(n35447), .Y(n26365) );
  AOI32XL U30556 ( .A0(n33788), .A1(n26367), .A2(n26366), .B0(conv_1[350]), 
        .B1(n26365), .Y(n26368) );
  NAND2XL U30557 ( .A(n26368), .B(n16652), .Y(n16113) );
  INVXL U30558 ( .A(conv_3[538]), .Y(n31284) );
  NAND2XL U30559 ( .A(conv_3[531]), .B(n26369), .Y(n27570) );
  NAND2XL U30560 ( .A(conv_3[533]), .B(n33718), .Y(n28960) );
  OAI2BB1XL U30561 ( .A0N(conv_3[535]), .A1N(n31142), .B0(n28959), .Y(n31185)
         );
  NAND4XL U30562 ( .A(conv_3[536]), .B(conv_3[537]), .C(n28959), .D(n31185), 
        .Y(n31286) );
  INVXL U30563 ( .A(conv_3[537]), .Y(n31171) );
  INVXL U30564 ( .A(conv_3[536]), .Y(n31190) );
  OAI21XL U30565 ( .A0(conv_3[535]), .A1(n31141), .B0(n33719), .Y(n31186) );
  NAND2XL U30566 ( .A(n31190), .B(n31186), .Y(n26370) );
  NAND2XL U30567 ( .A(n33719), .B(n26370), .Y(n31167) );
  NAND3XL U30568 ( .A(n33719), .B(n31171), .C(n31167), .Y(n31285) );
  NAND2XL U30569 ( .A(n31286), .B(n31285), .Y(n26372) );
  OAI21XL U30570 ( .A0(n16654), .A1(n26372), .B0(n31191), .Y(n26371) );
  AOI32XL U30571 ( .A0(n36020), .A1(n31284), .A2(n26372), .B0(conv_3[538]), 
        .B1(n26371), .Y(n26373) );
  NAND2XL U30572 ( .A(n26373), .B(n35588), .Y(n15385) );
  AOI22XL U30573 ( .A0(n36245), .A1(n34824), .B0(n34825), .B1(n26374), .Y(
        n34852) );
  INVXL U30574 ( .A(n34823), .Y(n26532) );
  NAND2XL U30575 ( .A(n34954), .B(n34847), .Y(n26530) );
  OAI211XL U30576 ( .A0(n34851), .A1(n28577), .B0(n26375), .C0(n26530), .Y(
        n26380) );
  INVXL U30577 ( .A(n34822), .Y(n34845) );
  AOI22XL U30578 ( .A0(n16665), .A1(n28406), .B0(n34984), .B1(n34845), .Y(
        n26378) );
  OAI21XL U30579 ( .A0(n35195), .A1(n26376), .B0(n34847), .Y(n26377) );
  OAI211XL U30580 ( .A0(n26531), .A1(n28479), .B0(n26378), .C0(n26377), .Y(
        n26379) );
  INVXL U30581 ( .A(n26541), .Y(n26389) );
  OAI2BB1XL U30582 ( .A0N(n28528), .A1N(n26538), .B0(n26383), .Y(n26388) );
  AOI222XL U30583 ( .A0(n26386), .A1(n36245), .B0(n26385), .B1(n22370), .C0(
        n26384), .C1(n28407), .Y(n26543) );
  OAI22XL U30584 ( .A0(n26543), .A1(n26575), .B0(n34989), .B1(n26542), .Y(
        n26387) );
  AOI32XL U30585 ( .A0(n22370), .A1(n28467), .A2(n26546), .B0(n26554), .B1(
        N18471), .Y(n26391) );
  AOI22XL U30586 ( .A0(n36245), .A1(n26393), .B0(n26392), .B1(n28292), .Y(
        n26394) );
  AOI21XL U30587 ( .A0(n22370), .A1(n26395), .B0(n26394), .Y(n26551) );
  OAI22XL U30588 ( .A0(n26551), .A1(n26575), .B0(n26550), .B1(n35135), .Y(
        n26396) );
  AOI222XL U30589 ( .A0(n26493), .A1(pool[11]), .B0(n26493), .B1(n34803), .C0(
        pool[11]), .C1(n34803), .Y(n26406) );
  OAI22XL U30590 ( .A0(n26401), .A1(n26474), .B0(n26400), .B1(n28479), .Y(
        n26403) );
  OAI22XL U30591 ( .A0(n26566), .A1(n26473), .B0(n26555), .B1(n28577), .Y(
        n26402) );
  AOI222XL U30592 ( .A0(n26406), .A1(n34804), .B0(n26406), .B1(n34805), .C0(
        n34804), .C1(n34805), .Y(n26407) );
  AOI222XL U30593 ( .A0(pool[13]), .A1(n28618), .B0(pool[13]), .B1(n26407), 
        .C0(n28618), .C1(n26407), .Y(n26461) );
  INVXL U30594 ( .A(n26574), .Y(n26416) );
  OAI21XL U30595 ( .A0(n26410), .A1(n26409), .B0(n26408), .Y(n26415) );
  AOI222XL U30596 ( .A0(n26413), .A1(n36245), .B0(n26412), .B1(n22370), .C0(
        n26411), .C1(n28407), .Y(n26576) );
  OAI22XL U30597 ( .A0(n26576), .A1(n26575), .B0(n26573), .B1(n35135), .Y(
        n26414) );
  OAI22XL U30598 ( .A0(n28489), .A1(n28577), .B0(n28491), .B1(n28553), .Y(
        n26420) );
  AOI2BB2XL U30599 ( .B0(n28494), .B1(n26451), .A0N(n26474), .A1N(n28488), .Y(
        n26418) );
  OAI211XL U30600 ( .A0(n28490), .A1(n26473), .B0(n26418), .C0(n26417), .Y(
        n26419) );
  AOI211XL U30601 ( .A0(n26470), .A1(n26421), .B0(n26420), .C0(n26419), .Y(
        n26438) );
  OAI22XL U30602 ( .A0(n28503), .A1(n28553), .B0(n26422), .B1(n28479), .Y(
        n26427) );
  AOI22XL U30603 ( .A0(n16667), .A1(n26587), .B0(n16671), .B1(n26423), .Y(
        n26425) );
  OAI211XL U30604 ( .A0(n28511), .A1(n34983), .B0(n26425), .C0(n26424), .Y(
        n26426) );
  OAI22XL U30605 ( .A0(n28469), .A1(n26474), .B0(n28472), .B1(n28577), .Y(
        n26431) );
  AOI22XL U30606 ( .A0(n28528), .A1(n28475), .B0(n16670), .B1(n28476), .Y(
        n26429) );
  OAI211XL U30607 ( .A0(n34989), .A1(n26582), .B0(n26429), .C0(n26428), .Y(
        n26430) );
  AOI211XL U30608 ( .A0(n34984), .A1(n26579), .B0(n26431), .C0(n26430), .Y(
        n26436) );
  AOI22XL U30609 ( .A0(n16667), .A1(n28437), .B0(n28436), .B1(n26451), .Y(
        n26435) );
  OAI22XL U30610 ( .A0(n28441), .A1(n26474), .B0(n28439), .B1(n26473), .Y(
        n26433) );
  OAI22XL U30611 ( .A0(n28440), .A1(n28479), .B0(n28449), .B1(n28553), .Y(
        n26432) );
  AOI211XL U30612 ( .A0(n26470), .A1(n26606), .B0(n26433), .C0(n26432), .Y(
        n26434) );
  OAI211XL U30613 ( .A0(n28438), .A1(n28575), .B0(n26435), .C0(n26434), .Y(
        n26484) );
  NAND4BXL U30614 ( .AN(n26484), .B(n26438), .C(n26437), .D(n26436), .Y(n26458) );
  AOI22XL U30615 ( .A0(n28528), .A1(n28514), .B0(n16671), .B1(n26439), .Y(
        n26443) );
  OAI22XL U30616 ( .A0(n28518), .A1(n26473), .B0(n28517), .B1(n34983), .Y(
        n26441) );
  OAI22XL U30617 ( .A0(n26610), .A1(n28575), .B0(n28519), .B1(n28577), .Y(
        n26440) );
  AOI211XL U30618 ( .A0(n16665), .A1(n28515), .B0(n26441), .C0(n26440), .Y(
        n26442) );
  OAI211XL U30619 ( .A0(n34989), .A1(n26615), .B0(n26443), .C0(n26442), .Y(
        n26483) );
  AOI22XL U30620 ( .A0(n34992), .A1(n28530), .B0(n26444), .B1(n26451), .Y(
        n26448) );
  OAI22XL U30621 ( .A0(n28531), .A1(n26474), .B0(n28532), .B1(n26473), .Y(
        n26446) );
  OAI2BB2XL U30622 ( .B0(n28533), .B1(n28577), .A0N(n28526), .A1N(n16670), .Y(
        n26445) );
  OAI211XL U30623 ( .A0(n34989), .A1(n26626), .B0(n26448), .C0(n26447), .Y(
        n26482) );
  AOI22XL U30624 ( .A0(n16667), .A1(n26450), .B0(n34984), .B1(n26449), .Y(
        n26456) );
  OAI2BB2XL U30625 ( .B0(n28457), .B1(n28575), .A0N(n28450), .A1N(n26451), .Y(
        n26454) );
  OAI22XL U30626 ( .A0(n26452), .A1(n28479), .B0(n28463), .B1(n28553), .Y(
        n26453) );
  AOI211XL U30627 ( .A0(n26470), .A1(n26618), .B0(n26454), .C0(n26453), .Y(
        n26455) );
  OAI211XL U30628 ( .A0(n28453), .A1(n26474), .B0(n26456), .C0(n26455), .Y(
        n26481) );
  NOR4BXL U30629 ( .AN(n28616), .B(n26483), .C(n26482), .D(n26481), .Y(n26457)
         );
  NAND2BXL U30630 ( .AN(n26458), .B(n26457), .Y(n26459) );
  AOI22XL U30631 ( .A0(n16667), .A1(n26632), .B0(n16670), .B1(n28410), .Y(
        n26466) );
  OAI22XL U30632 ( .A0(n28415), .A1(n26474), .B0(n34983), .B1(n26633), .Y(
        n26464) );
  OAI22XL U30633 ( .A0(n28417), .A1(n28479), .B0(n26462), .B1(n26473), .Y(
        n26463) );
  OAI211XL U30634 ( .A0(n34989), .A1(n26639), .B0(n26466), .C0(n26465), .Y(
        n26489) );
  INVXL U30635 ( .A(n26652), .Y(n26469) );
  OAI22XL U30636 ( .A0(n28550), .A1(n34983), .B0(n28554), .B1(n28577), .Y(
        n26468) );
  OAI22XL U30637 ( .A0(n28549), .A1(n26474), .B0(n28552), .B1(n28553), .Y(
        n26467) );
  AOI211XL U30638 ( .A0(n26470), .A1(n26469), .B0(n26468), .C0(n26467), .Y(
        n26471) );
  OAI211XL U30639 ( .A0(n28563), .A1(n26473), .B0(n26472), .C0(n26471), .Y(
        n26480) );
  AOI22XL U30640 ( .A0(n28528), .A1(n28573), .B0(n16670), .B1(n28574), .Y(
        n26478) );
  OAI22XL U30641 ( .A0(n26642), .A1(n34983), .B0(n28579), .B1(n28575), .Y(
        n26476) );
  OAI22XL U30642 ( .A0(n28580), .A1(n26474), .B0(n28576), .B1(n26473), .Y(
        n26475) );
  AOI211XL U30643 ( .A0(n28556), .A1(n28583), .B0(n26476), .C0(n26475), .Y(
        n26477) );
  OAI211XL U30644 ( .A0(n26479), .A1(n26647), .B0(n26478), .C0(n26477), .Y(
        n26485) );
  NOR3XL U30645 ( .A(pool[14]), .B(n26480), .C(n26485), .Y(n26488) );
  NAND4XL U30646 ( .A(pool[14]), .B(n26486), .C(n26485), .D(n26484), .Y(n26487) );
  NAND2XL U30647 ( .A(n34806), .B(pool[10]), .Y(n26492) );
  OAI21XL U30648 ( .A0(n26493), .A1(n34806), .B0(n26492), .Y(N29226) );
  AOI31XL U30649 ( .A0(conv_1[250]), .A1(conv_1[249]), .A2(n35411), .B0(n33663), .Y(n26971) );
  OAI21XL U30650 ( .A0(n26495), .A1(n36001), .B0(n35417), .Y(n26494) );
  NAND2XL U30651 ( .A(n26497), .B(n34682), .Y(n16212) );
  NAND2XL U30652 ( .A(n34721), .B(n27231), .Y(n26502) );
  NOR2X1 U30653 ( .A(n30195), .B(n33423), .Y(n27426) );
  NAND2XL U30654 ( .A(n27426), .B(conv_1[15]), .Y(n26498) );
  OR2XL U30655 ( .A(n26498), .B(n35272), .Y(n26500) );
  NAND2XL U30656 ( .A(n27429), .B(n26498), .Y(n26499) );
  NAND2XL U30657 ( .A(n27463), .B(conv_1[16]), .Y(n27462) );
  INVXL U30658 ( .A(conv_1[29]), .Y(n33443) );
  OAI21XL U30659 ( .A0(n26507), .A1(n16654), .B0(n35278), .Y(n26506) );
  NAND2XL U30660 ( .A(n26508), .B(n34544), .Y(n16443) );
  INVXL U30661 ( .A(conv_1[95]), .Y(n26777) );
  ADDFX1 U30662 ( .A(conv_1[93]), .B(n26511), .CI(n26510), .CO(n26512), .S(
        n22394) );
  OAI21XL U30663 ( .A0(n26517), .A1(n16655), .B0(n31361), .Y(n26516) );
  NAND2XL U30664 ( .A(n26518), .B(n34689), .Y(n16368) );
  AOI21XL U30665 ( .A0(n26520), .A1(n26519), .B0(n34775), .Y(n29286) );
  NOR2X1 U30666 ( .A(conv_1[414]), .B(n33385), .Y(n33386) );
  NAND2XL U30667 ( .A(conv_1[410]), .B(n26521), .Y(n29287) );
  NAND2XL U30668 ( .A(n35492), .B(conv_1[412]), .Y(n27596) );
  AOI21XL U30669 ( .A0(n33387), .A1(conv_1[414]), .B0(n35493), .Y(n29299) );
  AOI22XL U30670 ( .A0(n36020), .A1(n26522), .B0(conv_1[416]), .B1(n35495), 
        .Y(n26523) );
  NAND2XL U30671 ( .A(n26523), .B(n34689), .Y(n16047) );
  OAI21XL U30672 ( .A0(n26528), .A1(n16655), .B0(n35665), .Y(n26527) );
  NAND2XL U30673 ( .A(n26529), .B(n35588), .Y(n15603) );
  NAND2XL U30674 ( .A(n16721), .B(n34847), .Y(n34831) );
  OAI22XL U30675 ( .A0(n36245), .A1(n26530), .B0(n34831), .B1(n35135), .Y(
        n26536) );
  OAI22XL U30676 ( .A0(n34822), .A1(n28349), .B0(n34851), .B1(n28575), .Y(
        n26535) );
  OAI2BB2XL U30677 ( .B0(n26531), .B1(n28553), .A0N(n34846), .A1N(n28324), .Y(
        n26534) );
  AOI222XL U30678 ( .A0(n28406), .A1(n28291), .B0(n26532), .B1(n28290), .C0(
        n34847), .C1(n28289), .Y(n34853) );
  OAI22XL U30679 ( .A0(n34853), .A1(n28467), .B0(n26575), .B1(n34852), .Y(
        n26533) );
  AOI22XL U30680 ( .A0(n16665), .A1(n26538), .B0(n28324), .B1(n26537), .Y(
        n26540) );
  OAI211XL U30681 ( .A0(n26541), .A1(n34989), .B0(n26540), .C0(n26539), .Y(
        n26545) );
  OAI22XL U30682 ( .A0(n26543), .A1(n35159), .B0(n16701), .B1(n26542), .Y(
        n26544) );
  AOI22XL U30683 ( .A0(n16670), .A1(n26547), .B0(n28324), .B1(n26546), .Y(
        n26548) );
  OAI21XL U30684 ( .A0(n35135), .A1(n26549), .B0(n26548), .Y(n26553) );
  OAI22XL U30685 ( .A0(n26551), .A1(n35159), .B0(n26550), .B1(n34989), .Y(
        n26552) );
  AOI222XL U30686 ( .A0(pool[16]), .A1(n34807), .B0(pool[16]), .B1(n26666), 
        .C0(n34807), .C1(n26666), .Y(n26567) );
  OAI22XL U30687 ( .A0(n26556), .A1(n26621), .B0(n26555), .B1(n28575), .Y(
        n26560) );
  OAI22XL U30688 ( .A0(n26558), .A1(n28467), .B0(n26575), .B1(n26557), .Y(
        n26559) );
  NAND2XL U30689 ( .A(n16670), .B(n26563), .Y(n26564) );
  OAI211XL U30690 ( .A0(n26566), .A1(n28349), .B0(n26565), .C0(n26564), .Y(
        n34809) );
  AOI222XL U30691 ( .A0(n26567), .A1(n34809), .B0(n26567), .B1(n34811), .C0(
        n34809), .C1(n34811), .Y(n26568) );
  AOI222XL U30692 ( .A0(pool[18]), .A1(n27978), .B0(pool[18]), .B1(n26568), 
        .C0(n27978), .C1(n26568), .Y(n26631) );
  AOI22XL U30693 ( .A0(n16670), .A1(n26570), .B0(n28324), .B1(n26569), .Y(
        n26572) );
  OAI211XL U30694 ( .A0(n26573), .A1(n34989), .B0(n26572), .C0(n26571), .Y(
        n26578) );
  OAI22XL U30695 ( .A0(n26576), .A1(n35159), .B0(n26575), .B1(n26574), .Y(
        n26577) );
  OAI22XL U30696 ( .A0(n28469), .A1(n18196), .B0(n28472), .B1(n28575), .Y(
        n26584) );
  AOI22XL U30697 ( .A0(n16665), .A1(n28475), .B0(n18463), .B1(n28476), .Y(
        n26581) );
  AOI22XL U30698 ( .A0(n28366), .A1(n28473), .B0(n16663), .B1(n26579), .Y(
        n26580) );
  OAI211XL U30699 ( .A0(n26575), .A1(n26582), .B0(n26581), .C0(n26580), .Y(
        n26583) );
  AOI211XL U30700 ( .A0(n26585), .A1(n28372), .B0(n26584), .C0(n26583), .Y(
        n26603) );
  OAI22XL U30701 ( .A0(n28501), .A1(n18196), .B0(n28511), .B1(n28333), .Y(
        n26592) );
  AOI22XL U30702 ( .A0(n16670), .A1(n28498), .B0(n16663), .B1(n26588), .Y(
        n26589) );
  OAI211XL U30703 ( .A0(n28503), .A1(n16672), .B0(n26590), .C0(n26589), .Y(
        n26591) );
  AOI211XL U30704 ( .A0(n34827), .A1(n26593), .B0(n26592), .C0(n26591), .Y(
        n26602) );
  OAI22XL U30705 ( .A0(n28488), .A1(n18196), .B0(n28491), .B1(n16672), .Y(
        n26600) );
  AOI22XL U30706 ( .A0(n28366), .A1(n28486), .B0(n28494), .B1(n28372), .Y(
        n26597) );
  OAI211XL U30707 ( .A0(n26575), .A1(n26598), .B0(n26597), .C0(n26596), .Y(
        n26599) );
  AOI211XL U30708 ( .A0(n16665), .A1(n28487), .B0(n26600), .C0(n26599), .Y(
        n26601) );
  OAI22XL U30709 ( .A0(n28439), .A1(n28349), .B0(n28449), .B1(n16672), .Y(
        n26605) );
  OAI22XL U30710 ( .A0(n28438), .A1(n26621), .B0(n28440), .B1(n28553), .Y(
        n26604) );
  AOI211XL U30711 ( .A0(n34827), .A1(n26606), .B0(n26605), .C0(n26604), .Y(
        n26607) );
  OAI211XL U30712 ( .A0(n28441), .A1(n18196), .B0(n26608), .C0(n26607), .Y(
        n26658) );
  AOI22XL U30713 ( .A0(n16670), .A1(n28514), .B0(n26609), .B1(n28372), .Y(
        n26614) );
  OAI22XL U30714 ( .A0(n26610), .A1(n26621), .B0(n28519), .B1(n28575), .Y(
        n26612) );
  OAI22XL U30715 ( .A0(n28516), .A1(n18196), .B0(n28518), .B1(n28349), .Y(
        n26611) );
  AOI211XL U30716 ( .A0(n18463), .A1(n28515), .B0(n26612), .C0(n26611), .Y(
        n26613) );
  OAI211XL U30717 ( .A0(n26575), .A1(n26615), .B0(n26614), .C0(n26613), .Y(
        n26655) );
  AOI22XL U30718 ( .A0(n16670), .A1(n28451), .B0(n28450), .B1(n28372), .Y(
        n26620) );
  OAI22XL U30719 ( .A0(n28453), .A1(n18196), .B0(n28456), .B1(n28575), .Y(
        n26617) );
  OAI22XL U30720 ( .A0(n28455), .A1(n28349), .B0(n28463), .B1(n16672), .Y(
        n26616) );
  AOI211XL U30721 ( .A0(n34827), .A1(n26618), .B0(n26617), .C0(n26616), .Y(
        n26619) );
  OAI211XL U30722 ( .A0(n28457), .A1(n26621), .B0(n26620), .C0(n26619), .Y(
        n26653) );
  AOI22XL U30723 ( .A0(n16670), .A1(n28530), .B0(n28324), .B1(n28529), .Y(
        n26625) );
  OAI22XL U30724 ( .A0(n28532), .A1(n28349), .B0(n28531), .B1(n18196), .Y(
        n26623) );
  OAI22XL U30725 ( .A0(n28533), .A1(n28575), .B0(n28534), .B1(n28333), .Y(
        n26622) );
  AOI211XL U30726 ( .A0(n18463), .A1(n28526), .B0(n26623), .C0(n26622), .Y(
        n26624) );
  OAI211XL U30727 ( .A0(n26575), .A1(n26626), .B0(n26625), .C0(n26624), .Y(
        n26656) );
  NOR4XL U30728 ( .A(n26658), .B(n26655), .C(n26653), .D(n26656), .Y(n26627)
         );
  NAND2XL U30729 ( .A(n26628), .B(n26627), .Y(n26629) );
  OAI22XL U30730 ( .A0(n28417), .A1(n28553), .B0(n28333), .B1(n26633), .Y(
        n26636) );
  OAI22XL U30731 ( .A0(n28415), .A1(n18196), .B0(n26634), .B1(n16672), .Y(
        n26635) );
  AOI211XL U30732 ( .A0(n28366), .A1(n28412), .B0(n26636), .C0(n26635), .Y(
        n26637) );
  OAI211XL U30733 ( .A0(n26575), .A1(n26639), .B0(n26638), .C0(n26637), .Y(
        n26662) );
  AOI22XL U30734 ( .A0(n16670), .A1(n28573), .B0(n16663), .B1(n26640), .Y(
        n26646) );
  OAI22XL U30735 ( .A0(n26641), .A1(n16672), .B0(n28579), .B1(n26621), .Y(
        n26644) );
  OAI22XL U30736 ( .A0(n26642), .A1(n28333), .B0(n28580), .B1(n18196), .Y(
        n26643) );
  OAI211XL U30737 ( .A0(n26575), .A1(n26647), .B0(n26646), .C0(n26645), .Y(
        n26654) );
  AOI2BB2XL U30738 ( .B0(n28324), .B1(n28558), .A0N(n28349), .A1N(n28563), .Y(
        n26651) );
  OAI22XL U30739 ( .A0(n28550), .A1(n28333), .B0(n28554), .B1(n28575), .Y(
        n26649) );
  OAI22XL U30740 ( .A0(n28549), .A1(n18196), .B0(n28552), .B1(n16672), .Y(
        n26648) );
  AOI211XL U30741 ( .A0(n16665), .A1(n28560), .B0(n26649), .C0(n26648), .Y(
        n26650) );
  OAI211XL U30742 ( .A0(n16701), .A1(n26652), .B0(n26651), .C0(n26650), .Y(
        n26657) );
  NOR3XL U30743 ( .A(pool[19]), .B(n26654), .C(n26657), .Y(n26661) );
  NAND4XL U30744 ( .A(n26659), .B(n26658), .C(n26657), .D(n26656), .Y(n26660)
         );
  NAND2XL U30745 ( .A(n34810), .B(pool[15]), .Y(n26665) );
  OAI21XL U30746 ( .A0(n26666), .A1(n34810), .B0(n26665), .Y(N29231) );
  NAND3XL U30747 ( .A(conv_1[177]), .B(n26667), .C(n27538), .Y(n34685) );
  OR3XL U30748 ( .A(n26667), .B(conv_1[177]), .C(n27538), .Y(n34684) );
  INVXL U30749 ( .A(conv_1[178]), .Y(n34688) );
  AOI22XL U30750 ( .A0(conv_1[178]), .A1(n34685), .B0(n34684), .B1(n34688), 
        .Y(n26669) );
  NAND2XL U30751 ( .A(conv_1[179]), .B(n26669), .Y(n26668) );
  OAI211XL U30752 ( .A0(conv_1[179]), .A1(n26669), .B0(n33778), .C0(n26668), 
        .Y(n26670) );
  OAI211XL U30753 ( .A0(n34676), .A1(n26671), .B0(n34544), .C0(n26670), .Y(
        n16284) );
  INVXL U30754 ( .A(conv_1[235]), .Y(n26676) );
  NAND2XL U30755 ( .A(conv_1[235]), .B(n26674), .Y(n26673) );
  OAI211XL U30756 ( .A0(conv_1[235]), .A1(n26674), .B0(n33778), .C0(n26673), 
        .Y(n26675) );
  OAI211XL U30757 ( .A0(n35408), .A1(n26676), .B0(n34682), .C0(n26675), .Y(
        n16228) );
  INVXL U30758 ( .A(conv_3[521]), .Y(n26682) );
  NAND2XL U30759 ( .A(n31180), .B(n31292), .Y(n26678) );
  OAI21XL U30760 ( .A0(n31180), .A1(n31292), .B0(n26678), .Y(n26680) );
  AOI211XL U30761 ( .A0(n26682), .A1(n26680), .B0(n16654), .C0(n26679), .Y(
        n26681) );
  AOI2BB1XL U30762 ( .A0N(n26682), .A1N(n33303), .B0(n26681), .Y(n26683) );
  NAND2XL U30763 ( .A(n26683), .B(n35588), .Y(n15397) );
  INVXL U30764 ( .A(conv_1[92]), .Y(n26689) );
  NAND2XL U30765 ( .A(conv_1[92]), .B(n26687), .Y(n26686) );
  OAI211XL U30766 ( .A0(conv_1[92]), .A1(n26687), .B0(n33778), .C0(n26686), 
        .Y(n26688) );
  OAI211XL U30767 ( .A0(n31361), .A1(n26689), .B0(n26688), .C0(n33542), .Y(
        n16371) );
  INVXL U30768 ( .A(conv_1[150]), .Y(n26693) );
  OAI211XL U30769 ( .A0(conv_1[150]), .A1(n26691), .B0(n24499), .C0(n26690), 
        .Y(n26692) );
  OAI211XL U30770 ( .A0(n34048), .A1(n26693), .B0(n26692), .C0(n34773), .Y(
        n16313) );
  INVXL U30771 ( .A(conv_1[90]), .Y(n26697) );
  OAI211XL U30772 ( .A0(conv_1[90]), .A1(n26695), .B0(n16657), .C0(n26694), 
        .Y(n26696) );
  OAI211XL U30773 ( .A0(n31361), .A1(n26697), .B0(n26696), .C0(n34773), .Y(
        n16373) );
  INVXL U30774 ( .A(conv_1[91]), .Y(n26701) );
  OAI211XL U30775 ( .A0(conv_1[91]), .A1(n26699), .B0(n33778), .C0(n26698), 
        .Y(n26700) );
  OAI211XL U30776 ( .A0(n31361), .A1(n26701), .B0(n26700), .C0(n33067), .Y(
        n16372) );
  INVXL U30777 ( .A(n35022), .Y(n26706) );
  AOI22XL U30778 ( .A0(n35022), .A1(n26703), .B0(n26702), .B1(n26706), .Y(
        N29337) );
  AOI22XL U30779 ( .A0(n35022), .A1(n26705), .B0(n26704), .B1(n26706), .Y(
        N29339) );
  AOI22XL U30780 ( .A0(n35022), .A1(n26708), .B0(n26707), .B1(n26706), .Y(
        N29340) );
  NAND2BXL U30781 ( .AN(n26710), .B(n26709), .Y(n26712) );
  NAND2XL U30782 ( .A(n26714), .B(n26712), .Y(n26711) );
  OAI211XL U30783 ( .A0(n26714), .A1(n26712), .B0(n32656), .C0(n26711), .Y(
        n26713) );
  OAI211XL U30784 ( .A0(n34296), .A1(n26714), .B0(n16652), .C0(n26713), .Y(
        n16334) );
  INVXL U30785 ( .A(conv_3[349]), .Y(n26722) );
  AOI21XL U30786 ( .A0(n31391), .A1(n31392), .B0(n26718), .Y(n26720) );
  NAND2XL U30787 ( .A(conv_3[349]), .B(n26720), .Y(n26719) );
  OAI211XL U30788 ( .A0(conv_3[349]), .A1(n26720), .B0(n16656), .C0(n26719), 
        .Y(n26721) );
  OAI211XL U30789 ( .A0(n34746), .A1(n26722), .B0(n34097), .C0(n26721), .Y(
        n15756) );
  INVXL U30790 ( .A(conv_1[85]), .Y(n26728) );
  AOI21XL U30791 ( .A0(n26724), .A1(n34053), .B0(n26723), .Y(n26726) );
  NAND2XL U30792 ( .A(conv_1[85]), .B(n26726), .Y(n26725) );
  OAI211XL U30793 ( .A0(conv_1[85]), .A1(n26726), .B0(n32660), .C0(n26725), 
        .Y(n26727) );
  OAI211XL U30794 ( .A0(n34057), .A1(n26728), .B0(n34281), .C0(n26727), .Y(
        n16378) );
  INVXL U30795 ( .A(conv_1[86]), .Y(n26733) );
  NOR2BXL U30796 ( .AN(n26734), .B(n26729), .Y(n26731) );
  NAND2XL U30797 ( .A(conv_1[86]), .B(n26731), .Y(n26730) );
  OAI211XL U30798 ( .A0(conv_1[86]), .A1(n26731), .B0(n32181), .C0(n26730), 
        .Y(n26732) );
  OAI211XL U30799 ( .A0(n34057), .A1(n26733), .B0(n34544), .C0(n26732), .Y(
        n16377) );
  INVXL U30800 ( .A(conv_1[88]), .Y(n26832) );
  NAND4XL U30801 ( .A(conv_1[86]), .B(conv_1[87]), .C(n26735), .D(n26734), .Y(
        n26834) );
  NAND3XL U30802 ( .A(n26737), .B(n34053), .C(n26736), .Y(n26833) );
  NAND2XL U30803 ( .A(n26834), .B(n26833), .Y(n26739) );
  NAND2XL U30804 ( .A(conv_1[88]), .B(n26739), .Y(n26738) );
  OAI211XL U30805 ( .A0(conv_1[88]), .A1(n26739), .B0(n33822), .C0(n26738), 
        .Y(n26740) );
  OAI211XL U30806 ( .A0(n34057), .A1(n26832), .B0(n34281), .C0(n26740), .Y(
        n16375) );
  INVXL U30807 ( .A(conv_2[63]), .Y(n26747) );
  AOI21XL U30808 ( .A0(n26743), .A1(n26742), .B0(n26741), .Y(n26745) );
  NAND2XL U30809 ( .A(conv_2[63]), .B(n26745), .Y(n26744) );
  OAI211XL U30810 ( .A0(conv_2[63]), .A1(n26745), .B0(n24499), .C0(n26744), 
        .Y(n26746) );
  OAI211XL U30811 ( .A0(n35846), .A1(n26747), .B0(n34105), .C0(n26746), .Y(
        n15271) );
  INVXL U30812 ( .A(conv_1[138]), .Y(n26753) );
  XOR2XL U30813 ( .A(n26749), .B(n26748), .Y(n26751) );
  NAND2XL U30814 ( .A(conv_1[138]), .B(n26751), .Y(n26750) );
  OAI211XL U30815 ( .A0(conv_1[138]), .A1(n26751), .B0(n28751), .C0(n26750), 
        .Y(n26752) );
  OAI211XL U30816 ( .A0(n34271), .A1(n26753), .B0(n32867), .C0(n26752), .Y(
        n16325) );
  INVXL U30817 ( .A(conv_1[148]), .Y(n26825) );
  OAI2BB1XL U30818 ( .A0N(conv_1[145]), .A1N(n26754), .B0(n32780), .Y(n34266)
         );
  NAND4XL U30819 ( .A(conv_1[146]), .B(conv_1[147]), .C(n32780), .D(n34266), 
        .Y(n26827) );
  INVXL U30820 ( .A(conv_1[146]), .Y(n34272) );
  OAI21XL U30821 ( .A0(conv_1[145]), .A1(n26754), .B0(n35339), .Y(n34267) );
  AND2XL U30822 ( .A(n34272), .B(n34267), .Y(n26755) );
  NAND2XL U30823 ( .A(n35339), .B(n32781), .Y(n26826) );
  NAND2XL U30824 ( .A(n26827), .B(n26826), .Y(n26757) );
  NAND2XL U30825 ( .A(conv_1[148]), .B(n26757), .Y(n26756) );
  OAI211XL U30826 ( .A0(conv_1[148]), .A1(n26757), .B0(n33778), .C0(n26756), 
        .Y(n26758) );
  OAI211XL U30827 ( .A0(n34271), .A1(n26825), .B0(n34682), .C0(n26758), .Y(
        n16315) );
  AOI21XL U30828 ( .A0(n35339), .A1(n26760), .B0(n26759), .Y(n26762) );
  NAND2XL U30829 ( .A(conv_1[141]), .B(n26762), .Y(n26761) );
  OAI211XL U30830 ( .A0(conv_1[141]), .A1(n26762), .B0(n27932), .C0(n26761), 
        .Y(n26763) );
  OAI211XL U30831 ( .A0(n34271), .A1(n26764), .B0(n34696), .C0(n26763), .Y(
        n16322) );
  INVXL U30832 ( .A(conv_1[143]), .Y(n26770) );
  NAND2XL U30833 ( .A(conv_1[143]), .B(n26768), .Y(n26767) );
  OAI211XL U30834 ( .A0(conv_1[143]), .A1(n26768), .B0(n33822), .C0(n26767), 
        .Y(n26769) );
  OAI211XL U30835 ( .A0(n34271), .A1(n26770), .B0(n34544), .C0(n26769), .Y(
        n16320) );
  NAND2XL U30836 ( .A(n26772), .B(n26771), .Y(n26774) );
  NAND2XL U30837 ( .A(n26776), .B(n26774), .Y(n26773) );
  OAI211XL U30838 ( .A0(n26776), .A1(n26774), .B0(n34666), .C0(n26773), .Y(
        n26775) );
  OAI211XL U30839 ( .A0(n34271), .A1(n26776), .B0(n34682), .C0(n26775), .Y(
        n16323) );
  INVXL U30840 ( .A(conv_1[97]), .Y(n26812) );
  NAND2XL U30841 ( .A(conv_1[96]), .B(n26790), .Y(n26808) );
  NAND2XL U30842 ( .A(conv_1[98]), .B(n26784), .Y(n26795) );
  AOI21XL U30843 ( .A0(n31334), .A1(n26795), .B0(n26797), .Y(n26781) );
  NAND2XL U30844 ( .A(conv_1[99]), .B(n26781), .Y(n26780) );
  OAI211XL U30845 ( .A0(conv_1[99]), .A1(n26781), .B0(n33778), .C0(n26780), 
        .Y(n26782) );
  OAI211XL U30846 ( .A0(n31361), .A1(n26796), .B0(n34682), .C0(n26782), .Y(
        n16364) );
  AOI2BB1XL U30847 ( .A0N(n31337), .A1N(n26784), .B0(n26783), .Y(n26786) );
  NAND2XL U30848 ( .A(conv_1[98]), .B(n26786), .Y(n26785) );
  OAI211XL U30849 ( .A0(conv_1[98]), .A1(n26786), .B0(n24499), .C0(n26785), 
        .Y(n26787) );
  OAI211XL U30850 ( .A0(n31361), .A1(n26788), .B0(n34544), .C0(n26787), .Y(
        n16365) );
  INVXL U30851 ( .A(conv_1[96]), .Y(n26794) );
  AOI2BB1XL U30852 ( .A0N(n31337), .A1N(n26790), .B0(n26789), .Y(n26792) );
  NAND2XL U30853 ( .A(conv_1[96]), .B(n26792), .Y(n26791) );
  OAI211XL U30854 ( .A0(conv_1[96]), .A1(n26792), .B0(n28751), .C0(n26791), 
        .Y(n26793) );
  OAI211XL U30855 ( .A0(n31361), .A1(n26794), .B0(n16652), .C0(n26793), .Y(
        n16367) );
  AOI2BB1XL U30856 ( .A0N(n31337), .A1N(n26803), .B0(n26802), .Y(n26799) );
  NAND2XL U30857 ( .A(conv_1[100]), .B(n26799), .Y(n26798) );
  OAI211XL U30858 ( .A0(conv_1[100]), .A1(n26799), .B0(n30090), .C0(n26798), 
        .Y(n26800) );
  OAI211XL U30859 ( .A0(n31361), .A1(n26801), .B0(n34689), .C0(n26800), .Y(
        n16363) );
  INVXL U30860 ( .A(conv_1[101]), .Y(n26840) );
  OAI21XL U30861 ( .A0(conv_1[100]), .A1(n26802), .B0(n31337), .Y(n26839) );
  OAI2BB1XL U30862 ( .A0N(conv_1[100]), .A1N(n26803), .B0(n31334), .Y(n31333)
         );
  NAND2XL U30863 ( .A(n26839), .B(n31333), .Y(n26805) );
  NAND2XL U30864 ( .A(n26840), .B(n26805), .Y(n26804) );
  OAI211XL U30865 ( .A0(n26840), .A1(n26805), .B0(n33157), .C0(n26804), .Y(
        n26806) );
  OAI211XL U30866 ( .A0(n31361), .A1(n26840), .B0(n16652), .C0(n26806), .Y(
        n16362) );
  AOI21XL U30867 ( .A0(n31334), .A1(n26808), .B0(n26807), .Y(n26810) );
  NAND2XL U30868 ( .A(conv_1[97]), .B(n26810), .Y(n26809) );
  OAI211XL U30869 ( .A0(conv_1[97]), .A1(n26810), .B0(n33822), .C0(n26809), 
        .Y(n26811) );
  OAI211XL U30870 ( .A0(n31361), .A1(n26812), .B0(n34696), .C0(n26811), .Y(
        n16366) );
  INVXL U30871 ( .A(conv_3[409]), .Y(n26819) );
  AOI21XL U30872 ( .A0(n26815), .A1(n26814), .B0(n26813), .Y(n26817) );
  NAND2XL U30873 ( .A(conv_3[409]), .B(n26817), .Y(n26816) );
  OAI211XL U30874 ( .A0(conv_3[409]), .A1(n26817), .B0(n33778), .C0(n26816), 
        .Y(n26818) );
  OAI211XL U30875 ( .A0(n34227), .A1(n26819), .B0(n34097), .C0(n26818), .Y(
        n15752) );
  AOI21XL U30876 ( .A0(n35309), .A1(n27312), .B0(n26820), .Y(n26822) );
  NAND2XL U30877 ( .A(conv_1[52]), .B(n26822), .Y(n26821) );
  OAI211XL U30878 ( .A0(conv_1[52]), .A1(n26822), .B0(n32181), .C0(n26821), 
        .Y(n26823) );
  OAI211XL U30879 ( .A0(n35319), .A1(n26824), .B0(n34696), .C0(n26823), .Y(
        n16411) );
  AOI22XL U30880 ( .A0(conv_1[148]), .A1(n26827), .B0(n26826), .B1(n26825), 
        .Y(n26829) );
  NAND2XL U30881 ( .A(conv_1[149]), .B(n26829), .Y(n26828) );
  OAI211XL U30882 ( .A0(conv_1[149]), .A1(n26829), .B0(n32660), .C0(n26828), 
        .Y(n26830) );
  OAI211XL U30883 ( .A0(n34676), .A1(n26831), .B0(n34689), .C0(n26830), .Y(
        n16314) );
  AOI22XL U30884 ( .A0(conv_1[88]), .A1(n26834), .B0(n26833), .B1(n26832), .Y(
        n26836) );
  NAND2XL U30885 ( .A(conv_1[89]), .B(n26836), .Y(n26835) );
  OAI211XL U30886 ( .A0(conv_1[89]), .A1(n26836), .B0(n31735), .C0(n26835), 
        .Y(n26837) );
  OAI211XL U30887 ( .A0(n34676), .A1(n26838), .B0(n34281), .C0(n26837), .Y(
        n16374) );
  NAND2XL U30888 ( .A(n26840), .B(n26839), .Y(n26841) );
  AOI32XL U30889 ( .A0(conv_1[101]), .A1(n31335), .A2(n31333), .B0(n31337), 
        .B1(n31335), .Y(n26843) );
  AOI211XL U30890 ( .A0(n31336), .A1(n26843), .B0(n36042), .C0(n26842), .Y(
        n26844) );
  NAND2XL U30891 ( .A(n26845), .B(n34689), .Y(n16361) );
  NAND2X4 U30892 ( .A(n26852), .B(n26851), .Y(n26853) );
  OAI22XL U30893 ( .A0(n16645), .A1(n26854), .B0(n26867), .B1(n26910), .Y(
        n14585) );
  INVXL U30894 ( .A(weight_1[180]), .Y(n26863) );
  INVXL U30895 ( .A(weight_1[186]), .Y(n26865) );
  OAI22XL U30896 ( .A0(n16645), .A1(n26863), .B0(n26865), .B1(n26910), .Y(
        n14541) );
  INVXL U30897 ( .A(weight_1[240]), .Y(n26876) );
  INVXL U30898 ( .A(weight_1[246]), .Y(n26882) );
  OAI22XL U30899 ( .A0(n16650), .A1(n26876), .B0(n26882), .B1(n32777), .Y(
        n14551) );
  OAI22XL U30900 ( .A0(n16650), .A1(n26857), .B0(n26871), .B1(n26910), .Y(
        n14581) );
  OAI22XL U30901 ( .A0(n31084), .A1(n26885), .B0(n26854), .B1(n26910), .Y(
        n14584) );
  INVXL U30902 ( .A(weight_1[126]), .Y(n31318) );
  INVXL U30903 ( .A(weight_1[132]), .Y(n26855) );
  OAI22XL U30904 ( .A0(n16645), .A1(n31318), .B0(n26855), .B1(n16648), .Y(
        n14532) );
  INVXL U30905 ( .A(weight_1[258]), .Y(n26883) );
  INVXL U30906 ( .A(weight_1[264]), .Y(n26887) );
  OAI22XL U30907 ( .A0(n16650), .A1(n26883), .B0(n26887), .B1(n16647), .Y(
        n14554) );
  INVXL U30908 ( .A(weight_1[138]), .Y(n26856) );
  OAI22XL U30909 ( .A0(n16645), .A1(n26855), .B0(n26856), .B1(n16647), .Y(
        n14533) );
  INVXL U30910 ( .A(weight_1[144]), .Y(n26858) );
  OAI22XL U30911 ( .A0(n16645), .A1(n26856), .B0(n26858), .B1(n16647), .Y(
        n14534) );
  OAI22XL U30912 ( .A0(n16645), .A1(n26891), .B0(n26857), .B1(n26910), .Y(
        n14580) );
  INVXL U30913 ( .A(weight_1[150]), .Y(n26859) );
  OAI22XL U30914 ( .A0(n16645), .A1(n26858), .B0(n26859), .B1(n26910), .Y(
        n14535) );
  INVXL U30915 ( .A(weight_1[156]), .Y(n26860) );
  OAI22XL U30916 ( .A0(n16645), .A1(n26859), .B0(n26860), .B1(n32777), .Y(
        n14536) );
  INVXL U30917 ( .A(weight_1[162]), .Y(n26861) );
  OAI22XL U30918 ( .A0(n16645), .A1(n26860), .B0(n26861), .B1(n16648), .Y(
        n14537) );
  INVXL U30919 ( .A(weight_1[168]), .Y(n26862) );
  OAI22XL U30920 ( .A0(n16645), .A1(n26861), .B0(n26862), .B1(n32840), .Y(
        n14538) );
  INVXL U30921 ( .A(weight_1[174]), .Y(n26864) );
  OAI22XL U30922 ( .A0(n16645), .A1(n26862), .B0(n26864), .B1(n26910), .Y(
        n14539) );
  OAI22XL U30923 ( .A0(n16645), .A1(n26864), .B0(n26863), .B1(n26910), .Y(
        n14540) );
  INVXL U30924 ( .A(weight_1[378]), .Y(n26904) );
  INVXL U30925 ( .A(weight_1[384]), .Y(n26901) );
  OAI22XL U30926 ( .A0(n16650), .A1(n26904), .B0(n26901), .B1(n26910), .Y(
        n14574) );
  INVXL U30927 ( .A(weight_1[294]), .Y(n26878) );
  INVXL U30928 ( .A(weight_1[300]), .Y(n26903) );
  OAI22XL U30929 ( .A0(n32967), .A1(n26878), .B0(n26903), .B1(n26910), .Y(
        n14560) );
  OAI22XL U30930 ( .A0(n16645), .A1(n26865), .B0(n26868), .B1(n16648), .Y(
        n14542) );
  INVXL U30931 ( .A(weight_1[306]), .Y(n26902) );
  INVXL U30932 ( .A(weight_1[312]), .Y(n26866) );
  OAI22XL U30933 ( .A0(n16645), .A1(n26902), .B0(n26866), .B1(n32777), .Y(
        n14562) );
  INVXL U30934 ( .A(weight_1[318]), .Y(n26898) );
  OAI22XL U30935 ( .A0(n31077), .A1(n26866), .B0(n26898), .B1(n26910), .Y(
        n14563) );
  OAI22XL U30936 ( .A0(n16650), .A1(n26867), .B0(n26880), .B1(n26910), .Y(
        n14586) );
  INVXL U30937 ( .A(weight_1[462]), .Y(n26879) );
  OAI22XL U30938 ( .A0(n16645), .A1(n26879), .B0(n26907), .B1(n26910), .Y(
        n14588) );
  INVXL U30939 ( .A(weight_1[198]), .Y(n26869) );
  OAI22XL U30940 ( .A0(n16645), .A1(n26868), .B0(n26869), .B1(n26910), .Y(
        n14543) );
  INVXL U30941 ( .A(weight_1[204]), .Y(n26870) );
  OAI22XL U30942 ( .A0(n16650), .A1(n26869), .B0(n26870), .B1(n26910), .Y(
        n14544) );
  INVXL U30943 ( .A(weight_1[210]), .Y(n26872) );
  OAI22XL U30944 ( .A0(n16650), .A1(n26870), .B0(n26872), .B1(n16648), .Y(
        n14545) );
  OAI22XL U30945 ( .A0(n31071), .A1(n26871), .B0(n26886), .B1(n26910), .Y(
        n14582) );
  OAI22XL U30946 ( .A0(n16650), .A1(n26900), .B0(n26912), .B1(n26910), .Y(
        n14576) );
  INVXL U30947 ( .A(weight_1[216]), .Y(n26873) );
  OAI22XL U30948 ( .A0(n16650), .A1(n26872), .B0(n26873), .B1(n32840), .Y(
        n14546) );
  INVXL U30949 ( .A(weight_1[222]), .Y(n26874) );
  OAI22XL U30950 ( .A0(n16650), .A1(n26873), .B0(n26874), .B1(n26910), .Y(
        n14547) );
  INVXL U30951 ( .A(weight_1[228]), .Y(n26875) );
  OAI22XL U30952 ( .A0(n16650), .A1(n26874), .B0(n26875), .B1(n26910), .Y(
        n14548) );
  INVXL U30953 ( .A(weight_1[330]), .Y(n26889) );
  INVXL U30954 ( .A(weight_1[336]), .Y(n26894) );
  OAI22XL U30955 ( .A0(n31071), .A1(n26889), .B0(n26894), .B1(n26910), .Y(
        n14566) );
  INVXL U30956 ( .A(weight_1[342]), .Y(n26893) );
  INVXL U30957 ( .A(weight_1[348]), .Y(n26881) );
  OAI22XL U30958 ( .A0(n16650), .A1(n26893), .B0(n26881), .B1(n26910), .Y(
        n14568) );
  INVXL U30959 ( .A(weight_1[234]), .Y(n26877) );
  OAI22XL U30960 ( .A0(n16650), .A1(n26875), .B0(n26877), .B1(n16648), .Y(
        n14549) );
  OAI22XL U30961 ( .A0(n16650), .A1(n26877), .B0(n26876), .B1(n16647), .Y(
        n14550) );
  INVXL U30962 ( .A(weight_1[288]), .Y(n26895) );
  OAI22XL U30963 ( .A0(n31077), .A1(n26895), .B0(n26878), .B1(n32777), .Y(
        n14559) );
  OAI22XL U30964 ( .A0(n31084), .A1(n26880), .B0(n26879), .B1(n26910), .Y(
        n14587) );
  INVXL U30965 ( .A(weight_1[366]), .Y(n26908) );
  INVXL U30966 ( .A(weight_1[372]), .Y(n26905) );
  OAI22XL U30967 ( .A0(n16650), .A1(n26908), .B0(n26905), .B1(n26910), .Y(
        n14572) );
  INVXL U30968 ( .A(weight_1[354]), .Y(n26899) );
  OAI22XL U30969 ( .A0(n16650), .A1(n26881), .B0(n26899), .B1(n26910), .Y(
        n14569) );
  INVXL U30970 ( .A(weight_1[252]), .Y(n26884) );
  OAI22XL U30971 ( .A0(n16650), .A1(n26882), .B0(n26884), .B1(n16647), .Y(
        n14552) );
  OAI22XL U30972 ( .A0(n16650), .A1(n26884), .B0(n26883), .B1(n32777), .Y(
        n14553) );
  OAI22XL U30973 ( .A0(n16645), .A1(n26886), .B0(n26885), .B1(n26910), .Y(
        n14583) );
  INVXL U30974 ( .A(weight_1[270]), .Y(n26888) );
  OAI22XL U30975 ( .A0(n16650), .A1(n26887), .B0(n26888), .B1(n16647), .Y(
        n14555) );
  INVXL U30976 ( .A(weight_1[276]), .Y(n26890) );
  OAI22XL U30977 ( .A0(n32491), .A1(n26888), .B0(n26890), .B1(n16647), .Y(
        n14556) );
  INVXL U30978 ( .A(weight_1[324]), .Y(n26897) );
  OAI22XL U30979 ( .A0(n32491), .A1(n26897), .B0(n26889), .B1(n26910), .Y(
        n14565) );
  INVXL U30980 ( .A(weight_1[282]), .Y(n26896) );
  OAI22XL U30981 ( .A0(n31071), .A1(n26890), .B0(n26896), .B1(n16648), .Y(
        n14557) );
  OAI22XL U30982 ( .A0(n16650), .A1(n26911), .B0(n26892), .B1(n26910), .Y(
        n14578) );
  OAI22XL U30983 ( .A0(n16650), .A1(n26892), .B0(n26891), .B1(n26910), .Y(
        n14579) );
  OAI22XL U30984 ( .A0(n31077), .A1(n26894), .B0(n26893), .B1(n26910), .Y(
        n14567) );
  OAI22XL U30985 ( .A0(n26906), .A1(n26896), .B0(n26895), .B1(n16648), .Y(
        n14558) );
  OAI22XL U30986 ( .A0(n31071), .A1(n26898), .B0(n26897), .B1(n26910), .Y(
        n14564) );
  INVXL U30987 ( .A(weight_1[360]), .Y(n26909) );
  OAI22XL U30988 ( .A0(n16650), .A1(n26899), .B0(n26909), .B1(n26910), .Y(
        n14570) );
  OAI22XL U30989 ( .A0(n16650), .A1(n26901), .B0(n26900), .B1(n26910), .Y(
        n14575) );
  OAI22XL U30990 ( .A0(n31071), .A1(n26903), .B0(n26902), .B1(n32840), .Y(
        n14561) );
  OAI22XL U30991 ( .A0(n16650), .A1(n26905), .B0(n26904), .B1(n26910), .Y(
        n14573) );
  OAI22XL U30992 ( .A0(n31084), .A1(n26907), .B0(n26914), .B1(n16647), .Y(
        n14589) );
  OAI22XL U30993 ( .A0(n16650), .A1(n26909), .B0(n26908), .B1(n26910), .Y(
        n14571) );
  OAI22XL U30994 ( .A0(n16650), .A1(n26912), .B0(n26911), .B1(n26910), .Y(
        n14577) );
  OAI22XL U30995 ( .A0(n31071), .A1(n26913), .B0(n36124), .B1(n16647), .Y(
        n14591) );
  OAI22XL U30996 ( .A0(n16645), .A1(n26914), .B0(n16647), .B1(n26913), .Y(
        n14590) );
  INVXL U30997 ( .A(conv_1[137]), .Y(n26920) );
  NAND2XL U30998 ( .A(conv_1[137]), .B(n26918), .Y(n26917) );
  OAI211XL U30999 ( .A0(conv_1[137]), .A1(n26918), .B0(n32052), .C0(n26917), 
        .Y(n26919) );
  OAI211XL U31000 ( .A0(n34271), .A1(n26920), .B0(n33542), .C0(n26919), .Y(
        n16326) );
  INVXL U31001 ( .A(conv_1[94]), .Y(n26926) );
  NAND2XL U31002 ( .A(conv_1[94]), .B(n26924), .Y(n26923) );
  OAI211XL U31003 ( .A0(conv_1[94]), .A1(n26924), .B0(n33822), .C0(n26923), 
        .Y(n26925) );
  OAI211XL U31004 ( .A0(n31361), .A1(n26926), .B0(n35489), .C0(n26925), .Y(
        n16369) );
  INVXL U31005 ( .A(conv_1[139]), .Y(n26932) );
  NAND2XL U31006 ( .A(conv_1[139]), .B(n26930), .Y(n26929) );
  OAI211XL U31007 ( .A0(conv_1[139]), .A1(n26930), .B0(n32181), .C0(n26929), 
        .Y(n26931) );
  OAI211XL U31008 ( .A0(n34271), .A1(n26932), .B0(n35489), .C0(n26931), .Y(
        n16324) );
  INVXL U31009 ( .A(conv_2[227]), .Y(n26938) );
  NAND2XL U31010 ( .A(n26934), .B(n26933), .Y(n26936) );
  NAND2XL U31011 ( .A(n26938), .B(n26936), .Y(n26935) );
  OAI211XL U31012 ( .A0(n26938), .A1(n26936), .B0(n16657), .C0(n26935), .Y(
        n26937) );
  OAI211XL U31013 ( .A0(n34458), .A1(n26938), .B0(n34621), .C0(n26937), .Y(
        n15296) );
  INVXL U31014 ( .A(conv_1[438]), .Y(n26944) );
  NAND2XL U31015 ( .A(conv_1[438]), .B(n26942), .Y(n26941) );
  OAI211XL U31016 ( .A0(conv_1[438]), .A1(n26942), .B0(n28751), .C0(n26941), 
        .Y(n26943) );
  OAI211XL U31017 ( .A0(n35520), .A1(n26944), .B0(n26943), .C0(n32867), .Y(
        n16025) );
  NOR2BXL U31018 ( .AN(n26946), .B(n26945), .Y(n26948) );
  NAND2XL U31019 ( .A(conv_3[334]), .B(n26948), .Y(n26947) );
  OAI211XL U31020 ( .A0(conv_3[334]), .A1(n26948), .B0(n28751), .C0(n26947), 
        .Y(n26949) );
  OAI211XL U31021 ( .A0(n35748), .A1(n26950), .B0(n26949), .C0(n34097), .Y(
        n15757) );
  XOR2XL U31022 ( .A(n26952), .B(n26951), .Y(n26954) );
  NAND2XL U31023 ( .A(conv_1[468]), .B(n26954), .Y(n26953) );
  OAI211XL U31024 ( .A0(conv_1[468]), .A1(n26954), .B0(n28751), .C0(n26953), 
        .Y(n26955) );
  OAI211XL U31025 ( .A0(n33506), .A1(n26956), .B0(n26955), .C0(n32867), .Y(
        n15995) );
  NAND2XL U31026 ( .A(conv_1[0]), .B(n26957), .Y(n35271) );
  OAI211XL U31027 ( .A0(conv_1[0]), .A1(n26957), .B0(n33822), .C0(n35271), .Y(
        n26958) );
  OAI211XL U31028 ( .A0(n34552), .A1(n26959), .B0(n34773), .C0(n26958), .Y(
        n16463) );
  NAND3XL U31029 ( .A(conv_1[537]), .B(n26965), .C(n29236), .Y(n28001) );
  OR3XL U31030 ( .A(n26965), .B(conv_1[537]), .C(n29236), .Y(n28000) );
  NAND2XL U31031 ( .A(n28001), .B(n28000), .Y(n26962) );
  NAND2XL U31032 ( .A(conv_1[538]), .B(n26962), .Y(n26961) );
  OAI211XL U31033 ( .A0(conv_1[538]), .A1(n26962), .B0(n33788), .C0(n26961), 
        .Y(n26963) );
  OAI211XL U31034 ( .A0(n33432), .A1(n27999), .B0(n34696), .C0(n26963), .Y(
        n15925) );
  INVXL U31035 ( .A(conv_1[537]), .Y(n26969) );
  AOI21XL U31036 ( .A0(n26965), .A1(n29216), .B0(n26964), .Y(n26967) );
  NAND2XL U31037 ( .A(conv_1[537]), .B(n26967), .Y(n26966) );
  OAI211XL U31038 ( .A0(conv_1[537]), .A1(n26967), .B0(n27932), .C0(n26966), 
        .Y(n26968) );
  OAI211XL U31039 ( .A0(n33432), .A1(n26969), .B0(n16652), .C0(n26968), .Y(
        n15926) );
  NOR2X1 U31040 ( .A(n26972), .B(n26971), .Y(n33662) );
  NAND3XL U31041 ( .A(n33662), .B(conv_1[252]), .C(n35414), .Y(n27983) );
  NOR2X1 U31042 ( .A(n26972), .B(n35414), .Y(n33660) );
  NAND2XL U31043 ( .A(n33663), .B(n33661), .Y(n27982) );
  NAND2XL U31044 ( .A(n27983), .B(n27982), .Y(n26974) );
  OAI21XL U31045 ( .A0(n16655), .A1(n26974), .B0(n35417), .Y(n26973) );
  NAND2XL U31046 ( .A(n26975), .B(n34544), .Y(n16210) );
  INVXL U31047 ( .A(conv_1[33]), .Y(n26981) );
  XOR2XL U31048 ( .A(n26977), .B(n26976), .Y(n26979) );
  NAND2XL U31049 ( .A(conv_1[33]), .B(n26979), .Y(n26978) );
  OAI211XL U31050 ( .A0(conv_1[33]), .A1(n26979), .B0(n33822), .C0(n26978), 
        .Y(n26980) );
  OAI211XL U31051 ( .A0(n35302), .A1(n26981), .B0(n26980), .C0(n32867), .Y(
        n16430) );
  NAND2XL U31052 ( .A(conv_1[512]), .B(n26983), .Y(n26982) );
  OAI211XL U31053 ( .A0(conv_1[512]), .A1(n26983), .B0(n32181), .C0(n26982), 
        .Y(n26984) );
  OAI211XL U31054 ( .A0(n35547), .A1(n26985), .B0(n26984), .C0(n33542), .Y(
        n15951) );
  OAI211XL U31055 ( .A0(n26987), .A1(conv_1[467]), .B0(n28751), .C0(n26986), 
        .Y(n26988) );
  OAI211XL U31056 ( .A0(n33506), .A1(n26989), .B0(n26988), .C0(n33542), .Y(
        n15996) );
  INVXL U31057 ( .A(conv_1[62]), .Y(n26995) );
  NAND2XL U31058 ( .A(conv_1[62]), .B(n26993), .Y(n26992) );
  OAI211XL U31059 ( .A0(conv_1[62]), .A1(n26993), .B0(n31735), .C0(n26992), 
        .Y(n26994) );
  OAI211XL U31060 ( .A0(n35327), .A1(n26995), .B0(n26994), .C0(n33542), .Y(
        n16401) );
  INVXL U31061 ( .A(conv_1[77]), .Y(n26999) );
  NAND2XL U31062 ( .A(conv_1[77]), .B(n26997), .Y(n26996) );
  OAI211XL U31063 ( .A0(conv_1[77]), .A1(n26997), .B0(n33157), .C0(n26996), 
        .Y(n26998) );
  OAI211XL U31064 ( .A0(n34057), .A1(n26999), .B0(n26998), .C0(n33542), .Y(
        n16386) );
  INVXL U31065 ( .A(conv_1[439]), .Y(n27005) );
  NAND2XL U31066 ( .A(conv_1[439]), .B(n27003), .Y(n27002) );
  OAI211XL U31067 ( .A0(conv_1[439]), .A1(n27003), .B0(n28751), .C0(n27002), 
        .Y(n27004) );
  OAI211XL U31068 ( .A0(n35520), .A1(n27005), .B0(n27004), .C0(n35489), .Y(
        n16024) );
  NAND2XL U31069 ( .A(conv_1[469]), .B(n27009), .Y(n27008) );
  OAI211XL U31070 ( .A0(conv_1[469]), .A1(n27009), .B0(n28751), .C0(n27008), 
        .Y(n27010) );
  OAI211XL U31071 ( .A0(n33506), .A1(n27011), .B0(n27010), .C0(n35489), .Y(
        n15994) );
  OAI211XL U31072 ( .A0(n27013), .A1(conv_1[466]), .B0(n28751), .C0(n27012), 
        .Y(n27014) );
  OAI211XL U31073 ( .A0(n33506), .A1(n27015), .B0(n27014), .C0(n33067), .Y(
        n15997) );
  INVXL U31074 ( .A(conv_1[511]), .Y(n27019) );
  OAI211XL U31075 ( .A0(conv_1[511]), .A1(n27017), .B0(n33822), .C0(n27016), 
        .Y(n27018) );
  OAI211XL U31076 ( .A0(n35547), .A1(n27019), .B0(n27018), .C0(n33067), .Y(
        n15952) );
  INVXL U31077 ( .A(conv_1[61]), .Y(n27023) );
  OAI211XL U31078 ( .A0(conv_1[61]), .A1(n27021), .B0(n32611), .C0(n27020), 
        .Y(n27022) );
  OAI211XL U31079 ( .A0(n35327), .A1(n27023), .B0(n27022), .C0(n33067), .Y(
        n16402) );
  NAND2XL U31080 ( .A(n27025), .B(n27024), .Y(n27027) );
  NAND2XL U31081 ( .A(n27029), .B(n27027), .Y(n27026) );
  OAI211XL U31082 ( .A0(n27029), .A1(n27027), .B0(n32611), .C0(n27026), .Y(
        n27028) );
  OAI211XL U31083 ( .A0(n34057), .A1(n27029), .B0(n27028), .C0(n33067), .Y(
        n16387) );
  INVXL U31084 ( .A(conv_1[32]), .Y(n27035) );
  AND2XL U31085 ( .A(n27031), .B(n27030), .Y(n27033) );
  NAND2XL U31086 ( .A(conv_1[32]), .B(n27033), .Y(n27032) );
  OAI211XL U31087 ( .A0(conv_1[32]), .A1(n27033), .B0(n33778), .C0(n27032), 
        .Y(n27034) );
  OAI211XL U31088 ( .A0(n35302), .A1(n27035), .B0(n27034), .C0(n33542), .Y(
        n16431) );
  INVXL U31089 ( .A(conv_1[34]), .Y(n27041) );
  NAND2XL U31090 ( .A(conv_1[34]), .B(n27039), .Y(n27038) );
  OAI211XL U31091 ( .A0(conv_1[34]), .A1(n27039), .B0(n28751), .C0(n27038), 
        .Y(n27040) );
  OAI211XL U31092 ( .A0(n35302), .A1(n27041), .B0(n27040), .C0(n35489), .Y(
        n16429) );
  INVXL U31093 ( .A(conv_3[345]), .Y(n27045) );
  OAI211XL U31094 ( .A0(conv_3[345]), .A1(n27043), .B0(n33788), .C0(n27042), 
        .Y(n27044) );
  OAI211XL U31095 ( .A0(n34746), .A1(n27045), .B0(n27044), .C0(n34755), .Y(
        n15900) );
  NAND2XL U31096 ( .A(conv_2[257]), .B(n27047), .Y(n27046) );
  OAI211XL U31097 ( .A0(conv_2[257]), .A1(n27047), .B0(n33788), .C0(n27046), 
        .Y(n27048) );
  OAI211XL U31098 ( .A0(n34601), .A1(n27049), .B0(n27048), .C0(n34621), .Y(
        n15294) );
  INVXL U31099 ( .A(conv_2[212]), .Y(n27053) );
  NAND2XL U31100 ( .A(conv_2[212]), .B(n27051), .Y(n27050) );
  OAI211XL U31101 ( .A0(conv_2[212]), .A1(n27051), .B0(n33778), .C0(n27050), 
        .Y(n27052) );
  OAI211XL U31102 ( .A0(n35934), .A1(n27053), .B0(n27052), .C0(n34621), .Y(
        n15297) );
  NAND2XL U31103 ( .A(conv_2[527]), .B(n27055), .Y(n27054) );
  OAI211XL U31104 ( .A0(conv_2[527]), .A1(n27055), .B0(n32052), .C0(n27054), 
        .Y(n27056) );
  OAI211XL U31105 ( .A0(n34496), .A1(n27057), .B0(n27056), .C0(n34621), .Y(
        n15276) );
  INVXL U31106 ( .A(conv_3[300]), .Y(n27060) );
  OAI21XL U31107 ( .A0(n27058), .A1(n34389), .B0(n35736), .Y(n27059) );
  AOI32XL U31108 ( .A0(n33867), .A1(n27060), .A2(n34742), .B0(conv_3[300]), 
        .B1(n27059), .Y(n27061) );
  NAND2XL U31109 ( .A(n27061), .B(n34755), .Y(n15903) );
  INVXL U31110 ( .A(conv_3[510]), .Y(n27064) );
  OAI21XL U31111 ( .A0(n27062), .A1(n16655), .B0(n33303), .Y(n27063) );
  AOI32XL U31112 ( .A0(n34742), .A1(n27064), .A2(n34019), .B0(conv_3[510]), 
        .B1(n27063), .Y(n27065) );
  NAND2XL U31113 ( .A(n27065), .B(n34755), .Y(n15889) );
  AOI22XL U31114 ( .A0(n34948), .A1(n27067), .B0(n27066), .B1(n34945), .Y(
        N29310) );
  AOI22XL U31115 ( .A0(n34948), .A1(n27069), .B0(n27068), .B1(n34945), .Y(
        N29307) );
  INVXL U31116 ( .A(conv_1[5]), .Y(n27074) );
  AOI21XL U31117 ( .A0(intadd_2_n1), .A1(n27278), .B0(n27070), .Y(n27072) );
  NAND2XL U31118 ( .A(conv_1[5]), .B(n27072), .Y(n27071) );
  OAI211XL U31119 ( .A0(conv_1[5]), .A1(n27072), .B0(n32181), .C0(n27071), .Y(
        n27073) );
  OAI211XL U31120 ( .A0(n34552), .A1(n27074), .B0(n16652), .C0(n27073), .Y(
        n16458) );
  AOI2BB1XL U31121 ( .A0N(n27076), .A1N(n34547), .B0(n27075), .Y(n27078) );
  NAND2XL U31122 ( .A(conv_1[6]), .B(n27078), .Y(n27077) );
  OAI211XL U31123 ( .A0(conv_1[6]), .A1(n27078), .B0(n32181), .C0(n27077), .Y(
        n27079) );
  OAI211XL U31124 ( .A0(n34552), .A1(n27080), .B0(n34696), .C0(n27079), .Y(
        n16457) );
  INVXL U31125 ( .A(conv_2[183]), .Y(n27087) );
  ADDFXL U31126 ( .A(conv_2[182]), .B(n27082), .CI(n27081), .CO(n28651), .S(
        n23570) );
  AOI21XL U31127 ( .A0(n28651), .A1(n28652), .B0(n27083), .Y(n27085) );
  NAND2XL U31128 ( .A(conv_2[183]), .B(n27085), .Y(n27084) );
  OAI211XL U31129 ( .A0(conv_2[183]), .A1(n27085), .B0(n28751), .C0(n27084), 
        .Y(n27086) );
  OAI211XL U31130 ( .A0(n35917), .A1(n27087), .B0(n34105), .C0(n27086), .Y(
        n15263) );
  INVXL U31131 ( .A(conv_1[71]), .Y(n27093) );
  NAND2XL U31132 ( .A(conv_1[71]), .B(n27091), .Y(n27090) );
  OAI211XL U31133 ( .A0(conv_1[71]), .A1(n27091), .B0(n33157), .C0(n27090), 
        .Y(n27092) );
  OAI211XL U31134 ( .A0(n35327), .A1(n27093), .B0(n16652), .C0(n27092), .Y(
        n16392) );
  AOI21XL U31135 ( .A0(n35324), .A1(n27095), .B0(n27094), .Y(n27097) );
  NAND2XL U31136 ( .A(conv_1[69]), .B(n27097), .Y(n27096) );
  OAI211XL U31137 ( .A0(conv_1[69]), .A1(n27097), .B0(n33712), .C0(n27096), 
        .Y(n27098) );
  OAI211XL U31138 ( .A0(n35327), .A1(n27099), .B0(n34696), .C0(n27098), .Y(
        n16394) );
  AOI2BB1XL U31139 ( .A0N(n33638), .A1N(n27101), .B0(n27100), .Y(n27103) );
  NAND2XL U31140 ( .A(conv_1[66]), .B(n27103), .Y(n27102) );
  OAI211XL U31141 ( .A0(conv_1[66]), .A1(n27103), .B0(n32611), .C0(n27102), 
        .Y(n27104) );
  OAI211XL U31142 ( .A0(n35327), .A1(n27105), .B0(n34281), .C0(n27104), .Y(
        n16397) );
  NAND2XL U31143 ( .A(conv_1[65]), .B(n27109), .Y(n27108) );
  OAI211XL U31144 ( .A0(conv_1[65]), .A1(n27109), .B0(n33822), .C0(n27108), 
        .Y(n27110) );
  OAI211XL U31145 ( .A0(n35327), .A1(n27111), .B0(n16652), .C0(n27110), .Y(
        n16398) );
  NAND4XL U31146 ( .A(conv_1[506]), .B(conv_1[507]), .C(n27120), .D(n27132), 
        .Y(n27186) );
  INVXL U31147 ( .A(conv_1[507]), .Y(n27137) );
  NAND2XL U31148 ( .A(n27113), .B(n27112), .Y(n27114) );
  NAND3XL U31149 ( .A(n27131), .B(n27137), .C(n27133), .Y(n27185) );
  NAND2XL U31150 ( .A(n27186), .B(n27185), .Y(n27116) );
  NAND2XL U31151 ( .A(conv_1[508]), .B(n27116), .Y(n27115) );
  OAI211XL U31152 ( .A0(conv_1[508]), .A1(n27116), .B0(n33822), .C0(n27115), 
        .Y(n27117) );
  OAI211XL U31153 ( .A0(n33427), .A1(n27184), .B0(n16652), .C0(n27117), .Y(
        n15955) );
  OAI32XL U31154 ( .A0(n27120), .A1(conv_1[503]), .A2(n27119), .B0(n27131), 
        .B1(n27118), .Y(n27122) );
  NAND2XL U31155 ( .A(conv_1[504]), .B(n27122), .Y(n27121) );
  OAI211XL U31156 ( .A0(conv_1[504]), .A1(n27122), .B0(n33822), .C0(n27121), 
        .Y(n27123) );
  OAI211XL U31157 ( .A0(n33427), .A1(n27124), .B0(n16652), .C0(n27123), .Y(
        n15959) );
  OAI21XL U31158 ( .A0(n27131), .A1(n27126), .B0(n27125), .Y(n27128) );
  NAND2XL U31159 ( .A(n27130), .B(n27128), .Y(n27127) );
  OAI211XL U31160 ( .A0(n27130), .A1(n27128), .B0(n33822), .C0(n27127), .Y(
        n27129) );
  OAI211XL U31161 ( .A0(n33427), .A1(n27130), .B0(n34689), .C0(n27129), .Y(
        n15958) );
  AOI32XL U31162 ( .A0(conv_1[506]), .A1(n27133), .A2(n27132), .B0(n27131), 
        .B1(n27133), .Y(n27135) );
  NAND2XL U31163 ( .A(n27137), .B(n27135), .Y(n27134) );
  OAI211XL U31164 ( .A0(n27137), .A1(n27135), .B0(n33822), .C0(n27134), .Y(
        n27136) );
  OAI211XL U31165 ( .A0(n33427), .A1(n27137), .B0(n16652), .C0(n27136), .Y(
        n15956) );
  INVXL U31166 ( .A(conv_2[108]), .Y(n27144) );
  AOI21XL U31167 ( .A0(n27140), .A1(n27139), .B0(n27138), .Y(n27142) );
  NAND2XL U31168 ( .A(conv_2[108]), .B(n27142), .Y(n27141) );
  OAI211XL U31169 ( .A0(conv_2[108]), .A1(n27142), .B0(n32656), .C0(n27141), 
        .Y(n27143) );
  OAI211XL U31170 ( .A0(n35894), .A1(n27144), .B0(n34105), .C0(n27143), .Y(
        n15268) );
  INVXL U31171 ( .A(conv_1[447]), .Y(n27150) );
  INVXL U31172 ( .A(conv_1[444]), .Y(n27165) );
  OAI21XL U31173 ( .A0(conv_1[445]), .A1(n35513), .B0(n35515), .Y(n35521) );
  AOI32XL U31174 ( .A0(conv_1[446]), .A1(n27149), .A2(n35522), .B0(n35515), 
        .B1(n35523), .Y(n27147) );
  NAND2XL U31175 ( .A(n27150), .B(n27147), .Y(n27146) );
  OAI211XL U31176 ( .A0(n27150), .A1(n27147), .B0(n28751), .C0(n27146), .Y(
        n27148) );
  OAI211XL U31177 ( .A0(n35520), .A1(n27150), .B0(n16652), .C0(n27148), .Y(
        n16016) );
  INVXL U31178 ( .A(conv_1[448]), .Y(n27191) );
  NAND4XL U31179 ( .A(conv_1[446]), .B(conv_1[447]), .C(n27149), .D(n35522), 
        .Y(n27193) );
  NAND3XL U31180 ( .A(n35523), .B(n35515), .C(n27150), .Y(n27192) );
  NAND2XL U31181 ( .A(n27193), .B(n27192), .Y(n27152) );
  NAND2XL U31182 ( .A(conv_1[448]), .B(n27152), .Y(n27151) );
  OAI211XL U31183 ( .A0(conv_1[448]), .A1(n27152), .B0(n33822), .C0(n27151), 
        .Y(n27153) );
  OAI211XL U31184 ( .A0(n35520), .A1(n27191), .B0(n34544), .C0(n27153), .Y(
        n16015) );
  INVXL U31185 ( .A(conv_1[441]), .Y(n27159) );
  AOI2BB1XL U31186 ( .A0N(n35515), .A1N(n27155), .B0(n27154), .Y(n27157) );
  NAND2XL U31187 ( .A(conv_1[441]), .B(n27157), .Y(n27156) );
  OAI211XL U31188 ( .A0(conv_1[441]), .A1(n27157), .B0(n28751), .C0(n27156), 
        .Y(n27158) );
  OAI211XL U31189 ( .A0(n35520), .A1(n27159), .B0(n34544), .C0(n27158), .Y(
        n16022) );
  AOI21XL U31190 ( .A0(n27161), .A1(n35515), .B0(n27160), .Y(n27163) );
  NAND2XL U31191 ( .A(conv_1[444]), .B(n27163), .Y(n27162) );
  OAI211XL U31192 ( .A0(conv_1[444]), .A1(n27163), .B0(n28751), .C0(n27162), 
        .Y(n27164) );
  OAI211XL U31193 ( .A0(n35520), .A1(n27165), .B0(n34689), .C0(n27164), .Y(
        n16019) );
  NAND2XL U31194 ( .A(conv_1[440]), .B(n27169), .Y(n27168) );
  OAI211XL U31195 ( .A0(conv_1[440]), .A1(n27169), .B0(n28751), .C0(n27168), 
        .Y(n27170) );
  OAI211XL U31196 ( .A0(n35520), .A1(n27171), .B0(n34696), .C0(n27170), .Y(
        n16023) );
  AOI2BB1XL U31197 ( .A0N(n32887), .A1N(n27173), .B0(n27172), .Y(n27175) );
  NAND2XL U31198 ( .A(conv_1[473]), .B(n27175), .Y(n27174) );
  OAI211XL U31199 ( .A0(conv_1[473]), .A1(n27175), .B0(n32181), .C0(n27174), 
        .Y(n27176) );
  OAI211XL U31200 ( .A0(n33506), .A1(n27177), .B0(n16652), .C0(n27176), .Y(
        n15990) );
  AOI2BB1XL U31201 ( .A0N(n32887), .A1N(n27179), .B0(n27178), .Y(n27181) );
  NAND2XL U31202 ( .A(conv_1[471]), .B(n27181), .Y(n27180) );
  OAI211XL U31203 ( .A0(conv_1[471]), .A1(n27181), .B0(n28751), .C0(n27180), 
        .Y(n27182) );
  OAI211XL U31204 ( .A0(n33506), .A1(n27183), .B0(n16652), .C0(n27182), .Y(
        n15992) );
  AOI22XL U31205 ( .A0(conv_1[508]), .A1(n27186), .B0(n27185), .B1(n27184), 
        .Y(n27188) );
  NAND2XL U31206 ( .A(conv_1[509]), .B(n27188), .Y(n27187) );
  OAI211XL U31207 ( .A0(conv_1[509]), .A1(n27188), .B0(n33822), .C0(n27187), 
        .Y(n27189) );
  OAI211XL U31208 ( .A0(n33853), .A1(n27190), .B0(n34682), .C0(n27189), .Y(
        n15954) );
  AOI22XL U31209 ( .A0(conv_1[448]), .A1(n27193), .B0(n27192), .B1(n27191), 
        .Y(n27195) );
  NAND2XL U31210 ( .A(conv_1[449]), .B(n27195), .Y(n27194) );
  OAI211XL U31211 ( .A0(conv_1[449]), .A1(n27195), .B0(n33822), .C0(n27194), 
        .Y(n27196) );
  OAI211XL U31212 ( .A0(n33853), .A1(n27197), .B0(n16652), .C0(n27196), .Y(
        n16014) );
  AOI221XL U31213 ( .A0(n27199), .A1(n27932), .B0(n27198), .B1(n32660), .C0(
        n33633), .Y(n27204) );
  OAI211XL U31214 ( .A0(n33638), .A1(n27201), .B0(n32181), .C0(n27200), .Y(
        n27202) );
  OAI211XL U31215 ( .A0(n27204), .A1(n27203), .B0(n34696), .C0(n27202), .Y(
        n16395) );
  AOI22XL U31216 ( .A0(conv_1[73]), .A1(n27207), .B0(n27206), .B1(n27205), .Y(
        n27209) );
  NAND2XL U31217 ( .A(conv_1[74]), .B(n27209), .Y(n27208) );
  OAI211XL U31218 ( .A0(conv_1[74]), .A1(n27209), .B0(n32656), .C0(n27208), 
        .Y(n27210) );
  OAI211XL U31219 ( .A0(n34676), .A1(n27211), .B0(n34281), .C0(n27210), .Y(
        n16389) );
  INVXL U31220 ( .A(conv_1[485]), .Y(n29972) );
  OR2XL U31221 ( .A(n27212), .B(n27735), .Y(n33528) );
  OAI21XL U31222 ( .A0(n33403), .A1(n27735), .B0(n27215), .Y(n27216) );
  INVXL U31223 ( .A(n27216), .Y(n27374) );
  AOI222XL U31224 ( .A0(n27225), .A1(n27224), .B0(n27225), .B1(conv_1[483]), 
        .C0(n27224), .C1(conv_1[483]), .Y(n27217) );
  INVXL U31225 ( .A(n27217), .Y(n27218) );
  NOR2X1 U31226 ( .A(n27219), .B(n27218), .Y(n27399) );
  NAND2XL U31227 ( .A(conv_1[485]), .B(n27222), .Y(n27221) );
  OAI211XL U31228 ( .A0(conv_1[485]), .A1(n27222), .B0(n32181), .C0(n27221), 
        .Y(n27223) );
  OAI211XL U31229 ( .A0(n35544), .A1(n29972), .B0(n16652), .C0(n27223), .Y(
        n15978) );
  XOR2XL U31230 ( .A(n27225), .B(n27224), .Y(n27227) );
  NAND2XL U31231 ( .A(conv_1[483]), .B(n27227), .Y(n27226) );
  OAI211XL U31232 ( .A0(conv_1[483]), .A1(n27227), .B0(n32181), .C0(n27226), 
        .Y(n27228) );
  OAI211XL U31233 ( .A0(n35544), .A1(n27229), .B0(n32867), .C0(n27228), .Y(
        n15980) );
  NAND2XL U31234 ( .A(n27230), .B(n34444), .Y(n27237) );
  NAND2XL U31235 ( .A(n27231), .B(n34444), .Y(n27235) );
  NAND2XL U31236 ( .A(n27421), .B(n27429), .Y(n27232) );
  NAND2XL U31237 ( .A(n27435), .B(conv_1[451]), .Y(n27434) );
  AOI222XL U31238 ( .A0(n27380), .A1(conv_1[452]), .B0(n27380), .B1(n27379), 
        .C0(conv_1[452]), .C1(n27379), .Y(n27234) );
  NAND2XL U31239 ( .A(n27235), .B(n27234), .Y(n27250) );
  NOR2X1 U31240 ( .A(n27237), .B(n27236), .Y(n27392) );
  NAND2XL U31241 ( .A(n30048), .B(n30042), .Y(n30025) );
  NAND2XL U31242 ( .A(conv_1[456]), .B(n30019), .Y(n30050) );
  OAI21XL U31243 ( .A0(n28731), .A1(n30051), .B0(n28729), .Y(n27241) );
  NAND2XL U31244 ( .A(n28730), .B(n27241), .Y(n27240) );
  OAI211XL U31245 ( .A0(n28730), .A1(n27241), .B0(n28751), .C0(n27240), .Y(
        n27242) );
  OAI211XL U31246 ( .A0(n30056), .A1(n28730), .B0(n16652), .C0(n27242), .Y(
        n16001) );
  NAND2XL U31247 ( .A(conv_1[455]), .B(n27246), .Y(n27245) );
  OAI211XL U31248 ( .A0(conv_1[455]), .A1(n27246), .B0(n33822), .C0(n27245), 
        .Y(n27247) );
  OAI211XL U31249 ( .A0(n30056), .A1(n27248), .B0(n34682), .C0(n27247), .Y(
        n16008) );
  NOR2BXL U31250 ( .AN(n27250), .B(n27249), .Y(n27252) );
  NAND2XL U31251 ( .A(conv_1[453]), .B(n27252), .Y(n27251) );
  OAI211XL U31252 ( .A0(conv_1[453]), .A1(n27252), .B0(n33822), .C0(n27251), 
        .Y(n27253) );
  OAI211XL U31253 ( .A0(n30056), .A1(n27254), .B0(n32867), .C0(n27253), .Y(
        n16010) );
  AOI22XL U31254 ( .A0(n29246), .A1(conv_1[518]), .B0(n27259), .B1(n30267), 
        .Y(n27256) );
  NAND2XL U31255 ( .A(n27257), .B(n27256), .Y(n27255) );
  OAI211XL U31256 ( .A0(n27257), .A1(n27256), .B0(n32181), .C0(n27255), .Y(
        n27258) );
  OAI211XL U31257 ( .A0(n35547), .A1(n27259), .B0(n34544), .C0(n27258), .Y(
        n15945) );
  INVXL U31258 ( .A(conv_1[515]), .Y(n27265) );
  NAND2XL U31259 ( .A(conv_1[515]), .B(n27263), .Y(n27262) );
  OAI211XL U31260 ( .A0(conv_1[515]), .A1(n27263), .B0(n32181), .C0(n27262), 
        .Y(n27264) );
  OAI211XL U31261 ( .A0(n35547), .A1(n27265), .B0(n16652), .C0(n27264), .Y(
        n15948) );
  AOI2BB1XL U31262 ( .A0N(n29246), .A1N(n27267), .B0(n27266), .Y(n27269) );
  NAND2XL U31263 ( .A(conv_1[516]), .B(n27269), .Y(n27268) );
  OAI211XL U31264 ( .A0(conv_1[516]), .A1(n27269), .B0(n32181), .C0(n27268), 
        .Y(n27270) );
  OAI211XL U31265 ( .A0(n35547), .A1(n27271), .B0(n34689), .C0(n27270), .Y(
        n15947) );
  INVXL U31266 ( .A(conv_2[373]), .Y(n29466) );
  ADDFX1 U31267 ( .A(conv_2[370]), .B(n34570), .CI(n27272), .CO(n34571), .S(
        n23126) );
  NAND4XL U31268 ( .A(conv_2[371]), .B(conv_2[372]), .C(n34571), .D(n27273), 
        .Y(n29468) );
  NAND2XL U31269 ( .A(n29468), .B(n29467), .Y(n27275) );
  OAI21XL U31270 ( .A0(n16654), .A1(n27275), .B0(n36017), .Y(n27274) );
  AOI32XL U31271 ( .A0(n32052), .A1(n29466), .A2(n27275), .B0(conv_2[373]), 
        .B1(n27274), .Y(n27276) );
  NAND2XL U31272 ( .A(n27276), .B(n35859), .Y(n14955) );
  INVXL U31273 ( .A(conv_1[10]), .Y(n27283) );
  AOI21XL U31274 ( .A0(n27279), .A1(n27278), .B0(n27277), .Y(n27281) );
  NAND2XL U31275 ( .A(conv_1[10]), .B(n27281), .Y(n27280) );
  OAI211XL U31276 ( .A0(conv_1[10]), .A1(n27281), .B0(n33778), .C0(n27280), 
        .Y(n27282) );
  OAI211XL U31277 ( .A0(n34552), .A1(n27283), .B0(n34689), .C0(n27282), .Y(
        n16453) );
  INVXL U31278 ( .A(conv_1[7]), .Y(n27287) );
  NAND2XL U31279 ( .A(conv_1[7]), .B(n27285), .Y(n27284) );
  OAI211XL U31280 ( .A0(conv_1[7]), .A1(n27285), .B0(n33778), .C0(n27284), .Y(
        n27286) );
  OAI211XL U31281 ( .A0(n34552), .A1(n27287), .B0(n16652), .C0(n27286), .Y(
        n16456) );
  INVXL U31282 ( .A(conv_2[78]), .Y(n27293) );
  XOR2XL U31283 ( .A(n27289), .B(n27288), .Y(n27291) );
  NAND2XL U31284 ( .A(conv_2[78]), .B(n27291), .Y(n27290) );
  OAI211XL U31285 ( .A0(conv_2[78]), .A1(n27291), .B0(n33778), .C0(n27290), 
        .Y(n27292) );
  OAI211XL U31286 ( .A0(n35879), .A1(n27293), .B0(n34105), .C0(n27292), .Y(
        n15270) );
  NAND2XL U31287 ( .A(conv_1[35]), .B(n27297), .Y(n27296) );
  OAI211XL U31288 ( .A0(conv_1[35]), .A1(n27297), .B0(n33788), .C0(n27296), 
        .Y(n27298) );
  OAI211XL U31289 ( .A0(n35302), .A1(n27299), .B0(n34689), .C0(n27298), .Y(
        n16428) );
  AOI2BB1XL U31290 ( .A0N(n35296), .A1N(n27301), .B0(n27300), .Y(n27303) );
  NAND2XL U31291 ( .A(conv_1[38]), .B(n27303), .Y(n27302) );
  OAI211XL U31292 ( .A0(conv_1[38]), .A1(n27303), .B0(n27932), .C0(n27302), 
        .Y(n27304) );
  OAI211XL U31293 ( .A0(n35302), .A1(n27305), .B0(n34281), .C0(n27304), .Y(
        n16425) );
  AOI21XL U31294 ( .A0(n35289), .A1(n27307), .B0(n27306), .Y(n27309) );
  NAND2XL U31295 ( .A(conv_1[39]), .B(n27309), .Y(n27308) );
  OAI211XL U31296 ( .A0(conv_1[39]), .A1(n27309), .B0(n32181), .C0(n27308), 
        .Y(n27310) );
  OAI211XL U31297 ( .A0(n35302), .A1(n27311), .B0(n34689), .C0(n27310), .Y(
        n16424) );
  OAI211XL U31298 ( .A0(conv_1[51]), .A1(n27313), .B0(n30090), .C0(n27312), 
        .Y(n27314) );
  OAI211XL U31299 ( .A0(n35319), .A1(n27315), .B0(n34689), .C0(n27314), .Y(
        n16412) );
  AOI2BB1XL U31300 ( .A0N(n35316), .A1N(n27317), .B0(n27316), .Y(n27319) );
  NAND2XL U31301 ( .A(conv_1[53]), .B(n27319), .Y(n27318) );
  OAI211XL U31302 ( .A0(conv_1[53]), .A1(n27319), .B0(n32052), .C0(n27318), 
        .Y(n27320) );
  OAI211XL U31303 ( .A0(n35319), .A1(n27321), .B0(n34281), .C0(n27320), .Y(
        n16410) );
  OAI211XL U31304 ( .A0(conv_1[50]), .A1(n27323), .B0(n32181), .C0(n27322), 
        .Y(n27324) );
  OAI211XL U31305 ( .A0(n35319), .A1(n27325), .B0(n34544), .C0(n27324), .Y(
        n16413) );
  INVXL U31306 ( .A(conv_1[48]), .Y(n27331) );
  XOR2XL U31307 ( .A(n27327), .B(n27326), .Y(n27329) );
  NAND2XL U31308 ( .A(conv_1[48]), .B(n27329), .Y(n27328) );
  OAI211XL U31309 ( .A0(conv_1[48]), .A1(n27329), .B0(n34666), .C0(n27328), 
        .Y(n27330) );
  OAI211XL U31310 ( .A0(n35319), .A1(n27331), .B0(n32867), .C0(n27330), .Y(
        n16415) );
  NOR2X1 U31311 ( .A(n27608), .B(n30588), .Y(n35273) );
  INVXL U31312 ( .A(conv_1[22]), .Y(n27343) );
  NAND2XL U31313 ( .A(conv_1[21]), .B(n27345), .Y(n27339) );
  NAND2XL U31314 ( .A(conv_1[23]), .B(n27351), .Y(n27610) );
  AOI21XL U31315 ( .A0(conv_1[25]), .A1(n35274), .B0(n35275), .Y(n33202) );
  NAND2XL U31316 ( .A(conv_1[26]), .B(n27336), .Y(n27335) );
  OAI211XL U31317 ( .A0(conv_1[26]), .A1(n27336), .B0(n33778), .C0(n27335), 
        .Y(n27337) );
  OAI211XL U31318 ( .A0(n35278), .A1(n33201), .B0(n34281), .C0(n27337), .Y(
        n16437) );
  AOI21XL U31319 ( .A0(n30588), .A1(n27339), .B0(n27338), .Y(n27341) );
  NAND2XL U31320 ( .A(conv_1[22]), .B(n27341), .Y(n27340) );
  OAI211XL U31321 ( .A0(conv_1[22]), .A1(n27341), .B0(n33778), .C0(n27340), 
        .Y(n27342) );
  OAI211XL U31322 ( .A0(n35278), .A1(n27343), .B0(n16652), .C0(n27342), .Y(
        n16441) );
  AOI2BB1XL U31323 ( .A0N(n35275), .A1N(n27345), .B0(n27344), .Y(n27347) );
  NAND2XL U31324 ( .A(conv_1[21]), .B(n27347), .Y(n27346) );
  OAI211XL U31325 ( .A0(conv_1[21]), .A1(n27347), .B0(n33778), .C0(n27346), 
        .Y(n27348) );
  OAI211XL U31326 ( .A0(n35278), .A1(n27349), .B0(n34696), .C0(n27348), .Y(
        n16442) );
  AOI2BB1XL U31327 ( .A0N(n35275), .A1N(n27351), .B0(n27350), .Y(n27353) );
  NAND2XL U31328 ( .A(conv_1[23]), .B(n27353), .Y(n27352) );
  OAI211XL U31329 ( .A0(conv_1[23]), .A1(n27353), .B0(n33778), .C0(n27352), 
        .Y(n27354) );
  OAI211XL U31330 ( .A0(n35278), .A1(n27355), .B0(n34682), .C0(n27354), .Y(
        n16440) );
  INVXL U31331 ( .A(conv_1[18]), .Y(n27361) );
  NAND2XL U31332 ( .A(conv_1[18]), .B(n27359), .Y(n27358) );
  OAI211XL U31333 ( .A0(conv_1[18]), .A1(n27359), .B0(n33778), .C0(n27358), 
        .Y(n27360) );
  OAI211XL U31334 ( .A0(n35278), .A1(n27361), .B0(n32867), .C0(n27360), .Y(
        n16445) );
  AOI22XL U31335 ( .A0(conv_1[13]), .A1(n27364), .B0(n27363), .B1(n27362), .Y(
        n27366) );
  NAND2XL U31336 ( .A(conv_1[14]), .B(n27366), .Y(n27365) );
  OAI211XL U31337 ( .A0(conv_1[14]), .A1(n27366), .B0(n33778), .C0(n27365), 
        .Y(n27367) );
  OAI211XL U31338 ( .A0(n34676), .A1(n27368), .B0(n34682), .C0(n27367), .Y(
        n16449) );
  AOI22XL U31339 ( .A0(n34901), .A1(n27370), .B0(n27369), .B1(n34897), .Y(
        N29294) );
  AOI22XL U31340 ( .A0(n34901), .A1(n27372), .B0(n27371), .B1(n34897), .Y(
        N29295) );
  NAND2XL U31341 ( .A(conv_1[482]), .B(n27376), .Y(n27375) );
  OAI211XL U31342 ( .A0(conv_1[482]), .A1(n27376), .B0(n32181), .C0(n27375), 
        .Y(n27377) );
  OAI211XL U31343 ( .A0(n35544), .A1(n27378), .B0(n33542), .C0(n27377), .Y(
        n15981) );
  XOR2XL U31344 ( .A(n27380), .B(n27379), .Y(n27382) );
  NAND2XL U31345 ( .A(conv_1[452]), .B(n27382), .Y(n27381) );
  OAI211XL U31346 ( .A0(conv_1[452]), .A1(n27382), .B0(n33822), .C0(n27381), 
        .Y(n27383) );
  OAI211XL U31347 ( .A0(n30056), .A1(n27384), .B0(n33542), .C0(n27383), .Y(
        n16011) );
  AOI21XL U31348 ( .A0(n27387), .A1(n27386), .B0(n27385), .Y(n27389) );
  NAND2XL U31349 ( .A(conv_1[514]), .B(n27389), .Y(n27388) );
  OAI211XL U31350 ( .A0(conv_1[514]), .A1(n27389), .B0(n32181), .C0(n27388), 
        .Y(n27390) );
  OAI211XL U31351 ( .A0(n35547), .A1(n27391), .B0(n35489), .C0(n27390), .Y(
        n15949) );
  NAND2XL U31352 ( .A(conv_1[454]), .B(n27395), .Y(n27394) );
  OAI211XL U31353 ( .A0(conv_1[454]), .A1(n27395), .B0(n33822), .C0(n27394), 
        .Y(n27396) );
  OAI211XL U31354 ( .A0(n30056), .A1(n27397), .B0(n35489), .C0(n27396), .Y(
        n16009) );
  NAND2XL U31355 ( .A(conv_1[484]), .B(n27401), .Y(n27400) );
  OAI211XL U31356 ( .A0(conv_1[484]), .A1(n27401), .B0(n32181), .C0(n27400), 
        .Y(n27402) );
  OAI211XL U31357 ( .A0(n35544), .A1(n27403), .B0(n35489), .C0(n27402), .Y(
        n15979) );
  INVXL U31358 ( .A(conv_1[64]), .Y(n27410) );
  AOI21XL U31359 ( .A0(n27406), .A1(n27405), .B0(n27404), .Y(n27408) );
  NAND2XL U31360 ( .A(conv_1[64]), .B(n27408), .Y(n27407) );
  OAI211XL U31361 ( .A0(conv_1[64]), .A1(n27408), .B0(n32611), .C0(n27407), 
        .Y(n27409) );
  OAI211XL U31362 ( .A0(n35327), .A1(n27410), .B0(n35489), .C0(n27409), .Y(
        n16399) );
  INVXL U31363 ( .A(conv_2[287]), .Y(n27414) );
  OAI211XL U31364 ( .A0(n27412), .A1(conv_2[287]), .B0(n33822), .C0(n27411), 
        .Y(n27413) );
  OAI211XL U31365 ( .A0(n35963), .A1(n27414), .B0(n34621), .C0(n27413), .Y(
        n15292) );
  INVXL U31366 ( .A(conv_2[197]), .Y(n27420) );
  XOR2XL U31367 ( .A(n27416), .B(n27415), .Y(n27418) );
  NAND2XL U31368 ( .A(conv_2[197]), .B(n27418), .Y(n27417) );
  OAI211XL U31369 ( .A0(conv_2[197]), .A1(n27418), .B0(n32181), .C0(n27417), 
        .Y(n27419) );
  OAI211XL U31370 ( .A0(n35931), .A1(n27420), .B0(n34621), .C0(n27419), .Y(
        n15298) );
  OAI211XL U31371 ( .A0(n27422), .A1(conv_1[450]), .B0(n33822), .C0(n27421), 
        .Y(n27423) );
  OAI211XL U31372 ( .A0(n30056), .A1(n27424), .B0(n34773), .C0(n27423), .Y(
        n16013) );
  INVXL U31373 ( .A(conv_1[15]), .Y(n27427) );
  OAI21XL U31374 ( .A0(n16654), .A1(n27426), .B0(n35278), .Y(n27425) );
  NAND2XL U31375 ( .A(n27428), .B(n34773), .Y(n16448) );
  INVXL U31376 ( .A(n35271), .Y(n27430) );
  OAI32XL U31377 ( .A0(n35272), .A1(n27430), .A2(n35857), .B0(n35271), .B1(
        n27429), .Y(n35270) );
  NAND2XL U31378 ( .A(conv_1[1]), .B(n35270), .Y(n27431) );
  OAI211XL U31379 ( .A0(conv_1[1]), .A1(n35270), .B0(n32181), .C0(n27431), .Y(
        n27432) );
  OAI211XL U31380 ( .A0(n34552), .A1(n27433), .B0(n33067), .C0(n27432), .Y(
        n16462) );
  OAI211XL U31381 ( .A0(n27435), .A1(conv_1[451]), .B0(n33822), .C0(n27434), 
        .Y(n27436) );
  OAI211XL U31382 ( .A0(n30056), .A1(n27437), .B0(n33067), .C0(n27436), .Y(
        n16012) );
  INVXL U31383 ( .A(conv_1[47]), .Y(n27443) );
  NAND2XL U31384 ( .A(conv_1[47]), .B(n27441), .Y(n27440) );
  OAI211XL U31385 ( .A0(conv_1[47]), .A1(n27441), .B0(n34028), .C0(n27440), 
        .Y(n27442) );
  OAI211XL U31386 ( .A0(n35319), .A1(n27443), .B0(n33542), .C0(n27442), .Y(
        n16416) );
  INVXL U31387 ( .A(conv_1[17]), .Y(n27449) );
  XOR2XL U31388 ( .A(n27445), .B(n27444), .Y(n27447) );
  NAND2XL U31389 ( .A(conv_1[17]), .B(n27447), .Y(n27446) );
  OAI211XL U31390 ( .A0(conv_1[17]), .A1(n27447), .B0(n33778), .C0(n27446), 
        .Y(n27448) );
  OAI211XL U31391 ( .A0(n35278), .A1(n27449), .B0(n33542), .C0(n27448), .Y(
        n16446) );
  NAND2XL U31392 ( .A(conv_1[19]), .B(n27453), .Y(n27452) );
  OAI211XL U31393 ( .A0(conv_1[19]), .A1(n27453), .B0(n33778), .C0(n27452), 
        .Y(n27454) );
  OAI211XL U31394 ( .A0(n35278), .A1(n27455), .B0(n35489), .C0(n27454), .Y(
        n16444) );
  INVXL U31395 ( .A(conv_1[49]), .Y(n27461) );
  NAND2XL U31396 ( .A(conv_1[49]), .B(n27459), .Y(n27458) );
  OAI211XL U31397 ( .A0(conv_1[49]), .A1(n27459), .B0(n33788), .C0(n27458), 
        .Y(n27460) );
  OAI211XL U31398 ( .A0(n35319), .A1(n27461), .B0(n35489), .C0(n27460), .Y(
        n16414) );
  OAI211XL U31399 ( .A0(n27463), .A1(conv_1[16]), .B0(n33778), .C0(n27462), 
        .Y(n27464) );
  OAI211XL U31400 ( .A0(n35278), .A1(n27465), .B0(n33067), .C0(n27464), .Y(
        n16447) );
  NAND2XL U31401 ( .A(n27467), .B(n27466), .Y(n27469) );
  NAND2XL U31402 ( .A(n27471), .B(n27469), .Y(n27468) );
  OAI211XL U31403 ( .A0(n27471), .A1(n27469), .B0(n33982), .C0(n27468), .Y(
        n27470) );
  OAI211XL U31404 ( .A0(n35319), .A1(n27471), .B0(n33067), .C0(n27470), .Y(
        n16417) );
  AOI32XL U31405 ( .A0(n27474), .A1(n33427), .A2(n27472), .B0(n16654), .B1(
        n33427), .Y(n27476) );
  AOI22XL U31406 ( .A0(conv_1[497]), .A1(n27476), .B0(n27475), .B1(n27474), 
        .Y(n27477) );
  NAND2XL U31407 ( .A(n27477), .B(n33542), .Y(n15966) );
  NAND2XL U31408 ( .A(conv_3[166]), .B(n27481), .Y(n27480) );
  OAI211XL U31409 ( .A0(conv_3[166]), .A1(n27481), .B0(n34666), .C0(n27480), 
        .Y(n27482) );
  OAI211XL U31410 ( .A0(n35630), .A1(n27483), .B0(n27482), .C0(n33550), .Y(
        n15876) );
  INVXL U31411 ( .A(conv_3[181]), .Y(n27487) );
  NAND2XL U31412 ( .A(conv_3[181]), .B(n27485), .Y(n27484) );
  OAI211XL U31413 ( .A0(conv_3[181]), .A1(n27485), .B0(n27932), .C0(n27484), 
        .Y(n27486) );
  OAI211XL U31414 ( .A0(n34704), .A1(n27487), .B0(n27486), .C0(n33550), .Y(
        n15875) );
  INVXL U31415 ( .A(conv_3[61]), .Y(n27491) );
  NAND2XL U31416 ( .A(conv_3[61]), .B(n27489), .Y(n27488) );
  OAI211XL U31417 ( .A0(conv_3[61]), .A1(n27489), .B0(n33982), .C0(n27488), 
        .Y(n27490) );
  OAI211XL U31418 ( .A0(n35598), .A1(n27491), .B0(n27490), .C0(n33550), .Y(
        n15883) );
  INVXL U31419 ( .A(conv_3[210]), .Y(n27494) );
  OAI21XL U31420 ( .A0(n27492), .A1(n36042), .B0(n35665), .Y(n27493) );
  AOI32XL U31421 ( .A0(n34476), .A1(n27494), .A2(n34742), .B0(conv_3[210]), 
        .B1(n27493), .Y(n27495) );
  NAND2XL U31422 ( .A(n27495), .B(n34755), .Y(n15909) );
  INVXL U31423 ( .A(conv_3[151]), .Y(n27499) );
  OAI211XL U31424 ( .A0(n27497), .A1(conv_3[151]), .B0(n16656), .C0(n27496), 
        .Y(n27498) );
  OAI211XL U31425 ( .A0(n34751), .A1(n27499), .B0(n33550), .C0(n27498), .Y(
        n15877) );
  INVXL U31426 ( .A(conv_3[91]), .Y(n27503) );
  OAI211XL U31427 ( .A0(n27501), .A1(conv_3[91]), .B0(n32611), .C0(n27500), 
        .Y(n27502) );
  OAI211XL U31428 ( .A0(n35618), .A1(n27503), .B0(n33550), .C0(n27502), .Y(
        n15881) );
  INVXL U31429 ( .A(conv_3[196]), .Y(n27507) );
  OAI211XL U31430 ( .A0(n27505), .A1(conv_3[196]), .B0(n34028), .C0(n27504), 
        .Y(n27506) );
  OAI211XL U31431 ( .A0(n35646), .A1(n27507), .B0(n33550), .C0(n27506), .Y(
        n15874) );
  INVXL U31432 ( .A(conv_3[1]), .Y(n27512) );
  OAI211XL U31433 ( .A0(conv_3[1]), .A1(n27510), .B0(n33788), .C0(n27509), .Y(
        n27511) );
  OAI211XL U31434 ( .A0(n34383), .A1(n27512), .B0(n33550), .C0(n27511), .Y(
        n15887) );
  INVXL U31435 ( .A(conv_3[121]), .Y(n27518) );
  NOR2BXL U31436 ( .AN(n27514), .B(n27513), .Y(n27516) );
  NAND2XL U31437 ( .A(conv_3[121]), .B(n27516), .Y(n27515) );
  OAI211XL U31438 ( .A0(conv_3[121]), .A1(n27516), .B0(n16657), .C0(n27515), 
        .Y(n27517) );
  OAI211XL U31439 ( .A0(n35626), .A1(n27518), .B0(n33550), .C0(n27517), .Y(
        n15879) );
  INVXL U31440 ( .A(conv_3[106]), .Y(n27522) );
  OAI211XL U31441 ( .A0(n27520), .A1(conv_3[106]), .B0(n33788), .C0(n27519), 
        .Y(n27521) );
  OAI211XL U31442 ( .A0(n34200), .A1(n27522), .B0(n33550), .C0(n27521), .Y(
        n15880) );
  INVXL U31443 ( .A(conv_3[136]), .Y(n27526) );
  OAI211XL U31444 ( .A0(n27524), .A1(conv_3[136]), .B0(n34028), .C0(n27523), 
        .Y(n27525) );
  OAI211XL U31445 ( .A0(n34737), .A1(n27526), .B0(n33550), .C0(n27525), .Y(
        n15878) );
  INVXL U31446 ( .A(conv_3[31]), .Y(n27530) );
  OAI211XL U31447 ( .A0(n27528), .A1(conv_3[31]), .B0(n33712), .C0(n27527), 
        .Y(n27529) );
  OAI211XL U31448 ( .A0(n35594), .A1(n27530), .B0(n33550), .C0(n27529), .Y(
        n15885) );
  INVXL U31449 ( .A(conv_3[375]), .Y(n27536) );
  OAI21XL U31450 ( .A0(n27533), .A1(n16654), .B0(n34168), .Y(n27534) );
  AOI32XL U31451 ( .A0(n34742), .A1(n27536), .A2(n27535), .B0(conv_3[375]), 
        .B1(n27534), .Y(n27537) );
  NAND2XL U31452 ( .A(n27537), .B(n34755), .Y(n15898) );
  OAI2BB1XL U31453 ( .A0N(conv_1[172]), .A1N(n27539), .B0(n27538), .Y(n27541)
         );
  AOI31XL U31454 ( .A0(n36020), .A1(n27540), .A2(n27541), .B0(n35549), .Y(
        n27545) );
  OAI2BB1XL U31455 ( .A0N(n27542), .A1N(n27541), .B0(n28751), .Y(n27544) );
  AOI32XL U31456 ( .A0(n35346), .A1(n27545), .A2(n27544), .B0(n27543), .B1(
        n27545), .Y(n16290) );
  INVXL U31457 ( .A(conv_1[132]), .Y(n27548) );
  OAI21XL U31458 ( .A0(conv_1[131]), .A1(n30450), .B0(n34292), .Y(n27547) );
  INVXL U31459 ( .A(n34292), .Y(n30449) );
  OAI2BB1XL U31460 ( .A0N(conv_1[131]), .A1N(n30450), .B0(n30449), .Y(n27546)
         );
  AOI31XL U31461 ( .A0(n36020), .A1(n30451), .A2(n27546), .B0(n35549), .Y(
        n27550) );
  OAI2BB1XL U31462 ( .A0N(n27547), .A1N(n27546), .B0(n34028), .Y(n27549) );
  AOI32XL U31463 ( .A0(n34296), .A1(n27550), .A2(n27549), .B0(n27548), .B1(
        n27550), .Y(n16331) );
  NAND2XL U31464 ( .A(n33620), .B(n27555), .Y(n29076) );
  NAND2XL U31465 ( .A(n29080), .B(n29076), .Y(n29082) );
  OAI2BB1XL U31466 ( .A0N(conv_2[20]), .A1N(n29075), .B0(n28673), .Y(n29081)
         );
  NAND2XL U31467 ( .A(conv_2[21]), .B(n29081), .Y(n27831) );
  NAND2XL U31468 ( .A(n28673), .B(n27831), .Y(n27556) );
  AOI32XL U31469 ( .A0(n27831), .A1(n36020), .A2(n28673), .B0(n27557), .B1(
        n36020), .Y(n27558) );
  INVXL U31470 ( .A(conv_2[22]), .Y(n27832) );
  NOR2X1 U31471 ( .A(conv_1[262]), .B(n27564), .Y(n29197) );
  NAND2XL U31472 ( .A(n29203), .B(conv_1[261]), .Y(n29196) );
  NAND2XL U31473 ( .A(n29229), .B(n29196), .Y(n27563) );
  AOI32XL U31474 ( .A0(n29196), .A1(n36020), .A2(n29229), .B0(n27564), .B1(
        n36020), .Y(n27565) );
  AOI32XL U31475 ( .A0(n34080), .A1(n27566), .A2(n27565), .B0(n29195), .B1(
        n27566), .Y(n16201) );
  NAND2XL U31476 ( .A(n28959), .B(n27570), .Y(n27567) );
  AOI32XL U31477 ( .A0(n27570), .A1(n36020), .A2(n28959), .B0(n27569), .B1(
        n33712), .Y(n27572) );
  NAND2XL U31478 ( .A(n31363), .B(n27577), .Y(n27574) );
  AOI32XL U31479 ( .A0(n27577), .A1(n36020), .A2(n31363), .B0(n27576), .B1(
        n16657), .Y(n27579) );
  NAND2XL U31480 ( .A(n29328), .B(n27584), .Y(n27581) );
  AOI32XL U31481 ( .A0(n27584), .A1(n36020), .A2(n29328), .B0(n27583), .B1(
        n33157), .Y(n27586) );
  AOI32XL U31482 ( .A0(n35504), .A1(n27587), .A2(n27586), .B0(n27585), .B1(
        n27587), .Y(n16035) );
  ADDFXL U31483 ( .A(conv_3[337]), .B(n31980), .CI(n27588), .CO(n31962), .S(
        n23770) );
  NAND2XL U31484 ( .A(conv_3[338]), .B(n31962), .Y(n31956) );
  NAND2XL U31485 ( .A(n31967), .B(n31956), .Y(n27589) );
  AOI31XL U31486 ( .A0(n36020), .A1(n31955), .A2(n27589), .B0(n31384), .Y(
        n27592) );
  AOI32XL U31487 ( .A0(n31956), .A1(n36020), .A2(n31967), .B0(n27590), .B1(
        n36020), .Y(n27591) );
  NAND2XL U31488 ( .A(n34775), .B(n27596), .Y(n27593) );
  AOI31XL U31489 ( .A0(n36020), .A1(n27594), .A2(n27593), .B0(n35549), .Y(
        n27599) );
  AOI32XL U31490 ( .A0(n27596), .A1(n36020), .A2(n34775), .B0(n27595), .B1(
        n16656), .Y(n27598) );
  AOI32XL U31491 ( .A0(n35487), .A1(n27599), .A2(n27598), .B0(n27597), .B1(
        n27599), .Y(n16050) );
  NAND2XL U31492 ( .A(n29823), .B(n27603), .Y(n27600) );
  AOI31XL U31493 ( .A0(n36020), .A1(n27601), .A2(n27600), .B0(n35549), .Y(
        n27606) );
  AOI32XL U31494 ( .A0(n27603), .A1(n36020), .A2(n29823), .B0(n27602), .B1(
        n36020), .Y(n27605) );
  AOI32XL U31495 ( .A0(n33506), .A1(n27606), .A2(n27605), .B0(n27604), .B1(
        n27606), .Y(n15991) );
  NAND2XL U31496 ( .A(n30588), .B(n27610), .Y(n27607) );
  AOI31XL U31497 ( .A0(n36020), .A1(n27608), .A2(n27607), .B0(n35549), .Y(
        n27613) );
  AOI32XL U31498 ( .A0(n27610), .A1(n36020), .A2(n30588), .B0(n27609), .B1(
        n33712), .Y(n27612) );
  AOI32XL U31499 ( .A0(n35278), .A1(n27613), .A2(n27612), .B0(n27611), .B1(
        n27613), .Y(n16439) );
  INVXL U31500 ( .A(conv_3[488]), .Y(n33964) );
  ADDFXL U31501 ( .A(conv_3[485]), .B(n35831), .CI(n27614), .CO(n35822), .S(
        n23774) );
  OAI31XL U31502 ( .A0(conv_3[486]), .A1(conv_3[487]), .A2(n35822), .B0(n35831), .Y(n33959) );
  INVXL U31503 ( .A(n35831), .Y(n35823) );
  AOI21XL U31504 ( .A0(n33964), .A1(n33959), .B0(n35823), .Y(n27616) );
  NAND2XL U31505 ( .A(conv_3[486]), .B(n35817), .Y(n35821) );
  NAND2XL U31506 ( .A(conv_3[488]), .B(n33960), .Y(n31548) );
  NAND2XL U31507 ( .A(n35823), .B(n31548), .Y(n27615) );
  AOI31XL U31508 ( .A0(n36020), .A1(n31547), .A2(n27615), .B0(n16653), .Y(
        n27618) );
  AOI32XL U31509 ( .A0(n31548), .A1(n36020), .A2(n35823), .B0(n27616), .B1(
        n31735), .Y(n27617) );
  AOI32XL U31510 ( .A0(n35826), .A1(n27618), .A2(n27617), .B0(n31549), .B1(
        n27618), .Y(n15419) );
  INVXL U31511 ( .A(conv_3[509]), .Y(n34519) );
  NAND2XL U31512 ( .A(n29677), .B(n33424), .Y(n27624) );
  NAND2XL U31513 ( .A(n27619), .B(n33424), .Y(n27622) );
  NAND2XL U31514 ( .A(n31381), .B(conv_3[495]), .Y(n31380) );
  OAI21XL U31515 ( .A0(n30536), .A1(n33422), .B0(n31380), .Y(n30730) );
  NAND2XL U31516 ( .A(n27622), .B(n27621), .Y(n30724) );
  INVXL U31517 ( .A(conv_3[500]), .Y(n32075) );
  NAND2XL U31518 ( .A(conv_3[501]), .B(n35837), .Y(n32063) );
  NAND2XL U31519 ( .A(n33918), .B(n32063), .Y(n27628) );
  AOI31XL U31520 ( .A0(n36020), .A1(n32065), .A2(n27628), .B0(n16653), .Y(
        n27631) );
  AOI32XL U31521 ( .A0(n32063), .A1(n36020), .A2(n33918), .B0(n27629), .B1(
        n36020), .Y(n27630) );
  AOI32XL U31522 ( .A0(n35841), .A1(n27631), .A2(n27630), .B0(n32064), .B1(
        n27631), .Y(n15411) );
  NAND2XL U31523 ( .A(conv_1[396]), .B(n29269), .Y(n29356) );
  NAND2XL U31524 ( .A(n35471), .B(n29356), .Y(n27638) );
  AOI31XL U31525 ( .A0(n36020), .A1(n29358), .A2(n27638), .B0(n35549), .Y(
        n27641) );
  AOI32XL U31526 ( .A0(n29356), .A1(n36020), .A2(n35471), .B0(n27639), .B1(
        n16657), .Y(n27640) );
  INVXL U31527 ( .A(conv_1[397]), .Y(n29357) );
  AOI32XL U31528 ( .A0(n35477), .A1(n27641), .A2(n27640), .B0(n29357), .B1(
        n27641), .Y(n16066) );
  AOI21XL U31529 ( .A0(n30876), .A1(n33611), .B0(n27645), .Y(n27647) );
  NAND2XL U31530 ( .A(conv_2[455]), .B(n27647), .Y(n27646) );
  OAI211XL U31531 ( .A0(conv_2[455]), .A1(n27647), .B0(n16657), .C0(n27646), 
        .Y(n27648) );
  OAI211XL U31532 ( .A0(n34441), .A1(n27649), .B0(n34669), .C0(n27648), .Y(
        n14903) );
  NAND2XL U31533 ( .A(n30881), .B(n30877), .Y(n27666) );
  NAND2XL U31534 ( .A(n27676), .B(n27671), .Y(n27653) );
  AOI31XL U31535 ( .A0(conv_2[456]), .A1(conv_2[455]), .A2(n30876), .B0(n33611), .Y(n27665) );
  AOI21XL U31536 ( .A0(conv_2[458]), .A1(n27672), .B0(n33611), .Y(n27655) );
  AOI21XL U31537 ( .A0(n33611), .A1(n27653), .B0(n27655), .Y(n27651) );
  NAND2XL U31538 ( .A(conv_2[459]), .B(n27651), .Y(n27650) );
  OAI211XL U31539 ( .A0(conv_2[459]), .A1(n27651), .B0(n33712), .C0(n27650), 
        .Y(n27652) );
  OAI211XL U31540 ( .A0(n34441), .A1(n27654), .B0(n34669), .C0(n27652), .Y(
        n14899) );
  INVXL U31541 ( .A(n33611), .Y(n27677) );
  AOI21XL U31542 ( .A0(conv_2[460]), .A1(n33610), .B0(n33611), .Y(n27661) );
  NAND2XL U31543 ( .A(conv_2[461]), .B(n27657), .Y(n27656) );
  OAI211XL U31544 ( .A0(conv_2[461]), .A1(n27657), .B0(n32656), .C0(n27656), 
        .Y(n27658) );
  OAI211XL U31545 ( .A0(n34441), .A1(n27659), .B0(n34669), .C0(n27658), .Y(
        n14897) );
  AOI22XL U31546 ( .A0(n33611), .A1(n27680), .B0(n27678), .B1(n27677), .Y(
        n27663) );
  NAND2XL U31547 ( .A(n27679), .B(n27663), .Y(n27662) );
  OAI211XL U31548 ( .A0(n27679), .A1(n27663), .B0(n16657), .C0(n27662), .Y(
        n27664) );
  OAI211XL U31549 ( .A0(n34441), .A1(n27679), .B0(n34669), .C0(n27664), .Y(
        n14896) );
  AOI21XL U31550 ( .A0(n33611), .A1(n27666), .B0(n27665), .Y(n27668) );
  NAND2XL U31551 ( .A(conv_2[457]), .B(n27668), .Y(n27667) );
  OAI211XL U31552 ( .A0(conv_2[457]), .A1(n27668), .B0(n32660), .C0(n27667), 
        .Y(n27669) );
  OAI211XL U31553 ( .A0(n34441), .A1(n27670), .B0(n34669), .C0(n27669), .Y(
        n14901) );
  OAI21XL U31554 ( .A0(n33611), .A1(n27672), .B0(n27671), .Y(n27674) );
  NAND2XL U31555 ( .A(n27676), .B(n27674), .Y(n27673) );
  OAI211XL U31556 ( .A0(n27676), .A1(n27674), .B0(n34666), .C0(n27673), .Y(
        n27675) );
  OAI211XL U31557 ( .A0(n34441), .A1(n27676), .B0(n34669), .C0(n27675), .Y(
        n14900) );
  INVXL U31558 ( .A(conv_2[463]), .Y(n27958) );
  NAND3XL U31559 ( .A(n27678), .B(conv_2[462]), .C(n27677), .Y(n27960) );
  NAND3XL U31560 ( .A(n27680), .B(n33611), .C(n27679), .Y(n27959) );
  NAND2XL U31561 ( .A(n27960), .B(n27959), .Y(n27682) );
  NAND2XL U31562 ( .A(conv_2[463]), .B(n27682), .Y(n27681) );
  OAI211XL U31563 ( .A0(conv_2[463]), .A1(n27682), .B0(n32181), .C0(n27681), 
        .Y(n27683) );
  OAI211XL U31564 ( .A0(n34441), .A1(n27958), .B0(n34669), .C0(n27683), .Y(
        n14895) );
  AND2XL U31565 ( .A(n27687), .B(n27686), .Y(n28852) );
  INVXL U31566 ( .A(conv_2[534]), .Y(n29099) );
  INVXL U31567 ( .A(conv_2[532]), .Y(n29092) );
  NAND2XL U31568 ( .A(conv_2[531]), .B(n29625), .Y(n29088) );
  NAND2XL U31569 ( .A(conv_2[533]), .B(n33628), .Y(n29094) );
  AOI21XL U31570 ( .A0(conv_2[535]), .A1(n33373), .B0(n33629), .Y(n29100) );
  AOI22XL U31571 ( .A0(n33629), .A1(n28254), .B0(n28252), .B1(n29095), .Y(
        n27689) );
  NAND2XL U31572 ( .A(n28253), .B(n27689), .Y(n27688) );
  OAI211XL U31573 ( .A0(n28253), .A1(n27689), .B0(n27932), .C0(n27688), .Y(
        n27690) );
  OAI211XL U31574 ( .A0(n34496), .A1(n28253), .B0(n33815), .C0(n27690), .Y(
        n14846) );
  INVXL U31575 ( .A(conv_2[7]), .Y(n29587) );
  OAI31XL U31576 ( .A0(conv_2[5]), .A1(conv_2[6]), .A2(intadd_0_n1), .B0(
        n33571), .Y(n29581) );
  AOI21XL U31577 ( .A0(n29587), .A1(n29581), .B0(n29583), .Y(n33568) );
  AOI2BB1XL U31578 ( .A0N(conv_2[9]), .A1N(n28778), .B0(n29583), .Y(n28784) );
  OAI21XL U31579 ( .A0(conv_2[10]), .A1(n28784), .B0(n33571), .Y(n27695) );
  OAI2BB1XL U31580 ( .A0N(conv_2[5]), .A1N(intadd_0_n1), .B0(n29583), .Y(
        n28773) );
  NAND2XL U31581 ( .A(conv_2[6]), .B(n28773), .Y(n29582) );
  NAND2XL U31582 ( .A(conv_2[8]), .B(n33570), .Y(n28779) );
  OAI2BB1XL U31583 ( .A0N(conv_2[10]), .A1N(n28785), .B0(n29583), .Y(n29589)
         );
  NAND2XL U31584 ( .A(n27695), .B(n29589), .Y(n27693) );
  NAND2XL U31585 ( .A(n27696), .B(n27693), .Y(n27692) );
  OAI211XL U31586 ( .A0(n27696), .A1(n27693), .B0(n31735), .C0(n27692), .Y(
        n27694) );
  OAI211XL U31587 ( .A0(n30958), .A1(n27696), .B0(n33815), .C0(n27694), .Y(
        n15197) );
  NAND4XL U31588 ( .A(conv_2[11]), .B(conv_2[12]), .C(n29583), .D(n29589), .Y(
        n27930) );
  INVXL U31589 ( .A(conv_2[12]), .Y(n29594) );
  NAND2XL U31590 ( .A(n27696), .B(n27695), .Y(n27697) );
  NAND2XL U31591 ( .A(n33571), .B(n27697), .Y(n29590) );
  NAND3XL U31592 ( .A(n33571), .B(n29594), .C(n29590), .Y(n27929) );
  NAND2XL U31593 ( .A(n27930), .B(n27929), .Y(n27699) );
  NAND2XL U31594 ( .A(conv_2[13]), .B(n27699), .Y(n27698) );
  OAI211XL U31595 ( .A0(conv_2[13]), .A1(n27699), .B0(n31735), .C0(n27698), 
        .Y(n27700) );
  OAI211XL U31596 ( .A0(n30958), .A1(n27928), .B0(n35859), .C0(n27700), .Y(
        n15195) );
  INVXL U31597 ( .A(conv_2[42]), .Y(n27723) );
  INVXL U31598 ( .A(conv_2[37]), .Y(n27716) );
  INVXL U31599 ( .A(n27701), .Y(n27702) );
  OAI21XL U31600 ( .A0(n27704), .A1(n27703), .B0(n27702), .Y(n27705) );
  AND2XL U31601 ( .A(n27705), .B(n27706), .Y(n29701) );
  NAND2XL U31602 ( .A(conv_2[36]), .B(n27729), .Y(n27712) );
  NAND2XL U31603 ( .A(conv_2[38]), .B(n27718), .Y(n35861) );
  OAI2BB1XL U31604 ( .A0N(conv_2[40]), .A1N(n33587), .B0(n35862), .Y(n29617)
         );
  AOI32XL U31605 ( .A0(conv_2[41]), .A1(n35862), .A2(n29617), .B0(n33588), 
        .B1(n27724), .Y(n27709) );
  NAND2XL U31606 ( .A(n27723), .B(n27709), .Y(n27708) );
  OAI211XL U31607 ( .A0(n27723), .A1(n27709), .B0(n16657), .C0(n27708), .Y(
        n27710) );
  OAI211XL U31608 ( .A0(n35865), .A1(n27723), .B0(n34669), .C0(n27710), .Y(
        n15176) );
  AOI21XL U31609 ( .A0(n35862), .A1(n27712), .B0(n27711), .Y(n27714) );
  NAND2XL U31610 ( .A(conv_2[37]), .B(n27714), .Y(n27713) );
  OAI211XL U31611 ( .A0(conv_2[37]), .A1(n27714), .B0(n16657), .C0(n27713), 
        .Y(n27715) );
  OAI211XL U31612 ( .A0(n35865), .A1(n27716), .B0(n34669), .C0(n27715), .Y(
        n15181) );
  INVXL U31613 ( .A(conv_2[38]), .Y(n27722) );
  AOI2BB1XL U31614 ( .A0N(n33588), .A1N(n27718), .B0(n27717), .Y(n27720) );
  NAND2XL U31615 ( .A(conv_2[38]), .B(n27720), .Y(n27719) );
  OAI211XL U31616 ( .A0(conv_2[38]), .A1(n27720), .B0(n16657), .C0(n27719), 
        .Y(n27721) );
  OAI211XL U31617 ( .A0(n35865), .A1(n27722), .B0(n34669), .C0(n27721), .Y(
        n15180) );
  INVXL U31618 ( .A(conv_2[43]), .Y(n27951) );
  NAND4XL U31619 ( .A(conv_2[41]), .B(conv_2[42]), .C(n35862), .D(n29617), .Y(
        n27953) );
  NAND3XL U31620 ( .A(n27724), .B(n33588), .C(n27723), .Y(n27952) );
  NAND2XL U31621 ( .A(n27953), .B(n27952), .Y(n27726) );
  NAND2XL U31622 ( .A(conv_2[43]), .B(n27726), .Y(n27725) );
  OAI211XL U31623 ( .A0(conv_2[43]), .A1(n27726), .B0(n16657), .C0(n27725), 
        .Y(n27727) );
  OAI211XL U31624 ( .A0(n35865), .A1(n27951), .B0(n33815), .C0(n27727), .Y(
        n15175) );
  AOI2BB1XL U31625 ( .A0N(n33588), .A1N(n27729), .B0(n27728), .Y(n27731) );
  NAND2XL U31626 ( .A(conv_2[36]), .B(n27731), .Y(n27730) );
  OAI211XL U31627 ( .A0(conv_2[36]), .A1(n27731), .B0(n31735), .C0(n27730), 
        .Y(n27732) );
  OAI211XL U31628 ( .A0(n35865), .A1(n27733), .B0(n35859), .C0(n27732), .Y(
        n15182) );
  INVXL U31629 ( .A(conv_2[485]), .Y(n27746) );
  NAND2XL U31630 ( .A(n33530), .B(n28068), .Y(n27738) );
  OR2XL U31631 ( .A(n27734), .B(n18913), .Y(n30289) );
  OAI21XL U31632 ( .A0(n27735), .A1(n18913), .B0(n27734), .Y(n30288) );
  NAND2XL U31633 ( .A(conv_2[481]), .B(n30288), .Y(n27736) );
  AOI222XL U31634 ( .A0(n30338), .A1(conv_2[482]), .B0(n30338), .B1(n30337), 
        .C0(conv_2[482]), .C1(n30337), .Y(n27737) );
  NAND2XL U31635 ( .A(conv_2[485]), .B(n27743), .Y(n27742) );
  OAI211XL U31636 ( .A0(conv_2[485]), .A1(n27743), .B0(n16656), .C0(n27742), 
        .Y(n27744) );
  OAI211XL U31637 ( .A0(n34137), .A1(n27746), .B0(n34669), .C0(n27744), .Y(
        n14883) );
  AOI21XL U31638 ( .A0(conv_2[489]), .A1(n27753), .B0(n34132), .Y(n29577) );
  NAND2XL U31639 ( .A(conv_2[490]), .B(n27749), .Y(n27748) );
  OAI211XL U31640 ( .A0(conv_2[490]), .A1(n27749), .B0(n16656), .C0(n27748), 
        .Y(n27750) );
  OAI211XL U31641 ( .A0(n34137), .A1(n27751), .B0(n34669), .C0(n27750), .Y(
        n14878) );
  INVXL U31642 ( .A(conv_2[489]), .Y(n27757) );
  AOI21XL U31643 ( .A0(n27753), .A1(n34132), .B0(n27752), .Y(n27755) );
  NAND2XL U31644 ( .A(conv_2[489]), .B(n27755), .Y(n27754) );
  OAI211XL U31645 ( .A0(conv_2[489]), .A1(n27755), .B0(n16656), .C0(n27754), 
        .Y(n27756) );
  OAI211XL U31646 ( .A0(n34137), .A1(n27757), .B0(n34669), .C0(n27756), .Y(
        n14879) );
  INVXL U31647 ( .A(conv_2[487]), .Y(n27763) );
  NAND2XL U31648 ( .A(conv_2[487]), .B(n27761), .Y(n27760) );
  OAI211XL U31649 ( .A0(conv_2[487]), .A1(n27761), .B0(n16656), .C0(n27760), 
        .Y(n27762) );
  OAI211XL U31650 ( .A0(n34137), .A1(n27763), .B0(n34669), .C0(n27762), .Y(
        n14881) );
  INVXL U31651 ( .A(conv_2[521]), .Y(n31014) );
  INVXL U31652 ( .A(n27767), .Y(n27768) );
  NOR2X1 U31653 ( .A(conv_2[519]), .B(n28705), .Y(n28704) );
  OAI21XL U31654 ( .A0(conv_2[520]), .A1(n27793), .B0(n33580), .Y(n31009) );
  NAND2XL U31655 ( .A(n31014), .B(n31009), .Y(n27770) );
  INVXL U31656 ( .A(conv_2[519]), .Y(n28708) );
  INVXL U31657 ( .A(conv_2[517]), .Y(n27792) );
  INVXL U31658 ( .A(conv_2[515]), .Y(n27780) );
  NAND2XL U31659 ( .A(conv_2[516]), .B(n33579), .Y(n27788) );
  NAND2XL U31660 ( .A(conv_2[518]), .B(n27782), .Y(n28707) );
  OAI2BB1XL U31661 ( .A0N(conv_2[520]), .A1N(n27794), .B0(n28706), .Y(n31008)
         );
  AOI32XL U31662 ( .A0(conv_2[521]), .A1(n28202), .A2(n31008), .B0(n33580), 
        .B1(n28202), .Y(n27773) );
  NAND2XL U31663 ( .A(n28203), .B(n27773), .Y(n27772) );
  OAI211XL U31664 ( .A0(n28203), .A1(n27773), .B0(n16657), .C0(n27772), .Y(
        n27774) );
  OAI211XL U31665 ( .A0(n31013), .A1(n28203), .B0(n34669), .C0(n27774), .Y(
        n14856) );
  NAND2XL U31666 ( .A(conv_2[515]), .B(n27778), .Y(n27777) );
  OAI211XL U31667 ( .A0(conv_2[515]), .A1(n27778), .B0(n33822), .C0(n27777), 
        .Y(n27779) );
  OAI211XL U31668 ( .A0(n31013), .A1(n27780), .B0(n34669), .C0(n27779), .Y(
        n14863) );
  INVXL U31669 ( .A(conv_2[518]), .Y(n27786) );
  AOI2BB1XL U31670 ( .A0N(n33580), .A1N(n27782), .B0(n27781), .Y(n27784) );
  NAND2XL U31671 ( .A(conv_2[518]), .B(n27784), .Y(n27783) );
  OAI211XL U31672 ( .A0(conv_2[518]), .A1(n27784), .B0(n32611), .C0(n27783), 
        .Y(n27785) );
  OAI211XL U31673 ( .A0(n31013), .A1(n27786), .B0(n34669), .C0(n27785), .Y(
        n14860) );
  AOI21XL U31674 ( .A0(n28706), .A1(n27788), .B0(n27787), .Y(n27790) );
  NAND2XL U31675 ( .A(conv_2[517]), .B(n27790), .Y(n27789) );
  OAI211XL U31676 ( .A0(conv_2[517]), .A1(n27790), .B0(n34028), .C0(n27789), 
        .Y(n27791) );
  OAI211XL U31677 ( .A0(n31013), .A1(n27792), .B0(n34669), .C0(n27791), .Y(
        n14861) );
  NAND2XL U31678 ( .A(conv_2[520]), .B(n27796), .Y(n27795) );
  OAI211XL U31679 ( .A0(conv_2[520]), .A1(n27796), .B0(n16657), .C0(n27795), 
        .Y(n27797) );
  OAI211XL U31680 ( .A0(n31013), .A1(n27798), .B0(n34669), .C0(n27797), .Y(
        n14858) );
  AOI222XL U31681 ( .A0(conv_2[49]), .A1(n29739), .B0(conv_2[49]), .B1(n29740), 
        .C0(n29739), .C1(n29740), .Y(n27802) );
  NOR2X1 U31682 ( .A(n31134), .B(n27802), .Y(n27806) );
  NAND2XL U31683 ( .A(conv_2[50]), .B(n27804), .Y(n27803) );
  OAI211XL U31684 ( .A0(conv_2[50]), .A1(n27804), .B0(n16657), .C0(n27803), 
        .Y(n27805) );
  OAI211XL U31685 ( .A0(n34505), .A1(n27808), .B0(n34669), .C0(n27805), .Y(
        n15173) );
  INVXL U31686 ( .A(conv_2[55]), .Y(n27812) );
  AOI2BB1XL U31687 ( .A0N(n27808), .A1N(n27807), .B0(n31137), .Y(n27820) );
  NAND2XL U31688 ( .A(conv_2[53]), .B(n27814), .Y(n28714) );
  NOR2X1 U31689 ( .A(n28712), .B(n31134), .Y(n27825) );
  AOI2BB1XL U31690 ( .A0N(n31137), .A1N(n27826), .B0(n27825), .Y(n27810) );
  NAND2XL U31691 ( .A(conv_2[55]), .B(n27810), .Y(n27809) );
  OAI211XL U31692 ( .A0(conv_2[55]), .A1(n27810), .B0(n16657), .C0(n27809), 
        .Y(n27811) );
  OAI211XL U31693 ( .A0(n34505), .A1(n27812), .B0(n33815), .C0(n27811), .Y(
        n15168) );
  INVXL U31694 ( .A(conv_2[53]), .Y(n27818) );
  AOI21XL U31695 ( .A0(n27814), .A1(n31137), .B0(n27813), .Y(n27816) );
  NAND2XL U31696 ( .A(conv_2[53]), .B(n27816), .Y(n27815) );
  OAI211XL U31697 ( .A0(conv_2[53]), .A1(n27816), .B0(n16657), .C0(n27815), 
        .Y(n27817) );
  OAI211XL U31698 ( .A0(n34505), .A1(n27818), .B0(n35859), .C0(n27817), .Y(
        n15170) );
  NAND2XL U31699 ( .A(conv_2[51]), .B(n27822), .Y(n27821) );
  OAI211XL U31700 ( .A0(conv_2[51]), .A1(n27822), .B0(n16657), .C0(n27821), 
        .Y(n27823) );
  OAI211XL U31701 ( .A0(n34505), .A1(n27824), .B0(n33815), .C0(n27823), .Y(
        n15172) );
  OAI21XL U31702 ( .A0(conv_2[55]), .A1(n27825), .B0(n31137), .Y(n30160) );
  OAI2BB1XL U31703 ( .A0N(conv_2[55]), .A1N(n27826), .B0(n31134), .Y(n31133)
         );
  NAND2XL U31704 ( .A(n30160), .B(n31133), .Y(n27828) );
  NAND2XL U31705 ( .A(n30161), .B(n27828), .Y(n27827) );
  OAI211XL U31706 ( .A0(n30161), .A1(n27828), .B0(n16657), .C0(n27827), .Y(
        n27829) );
  OAI211XL U31707 ( .A0(n34505), .A1(n30161), .B0(n34735), .C0(n27829), .Y(
        n15167) );
  INVXL U31708 ( .A(conv_2[28]), .Y(n27936) );
  NAND2XL U31709 ( .A(conv_2[23]), .B(n33619), .Y(n28674) );
  AOI21XL U31710 ( .A0(conv_2[25]), .A1(n27917), .B0(n33620), .Y(n27836) );
  NAND3XL U31711 ( .A(n27842), .B(conv_2[27]), .C(n28673), .Y(n27938) );
  INVXL U31712 ( .A(conv_2[27]), .Y(n27847) );
  NAND3XL U31713 ( .A(n27843), .B(n33620), .C(n27847), .Y(n27937) );
  NAND2XL U31714 ( .A(n27938), .B(n27937), .Y(n27834) );
  NAND2XL U31715 ( .A(conv_2[28]), .B(n27834), .Y(n27833) );
  OAI211XL U31716 ( .A0(conv_2[28]), .A1(n27834), .B0(n16656), .C0(n27833), 
        .Y(n27835) );
  OAI211XL U31717 ( .A0(n30412), .A1(n27936), .B0(n34669), .C0(n27835), .Y(
        n15185) );
  NAND2XL U31718 ( .A(conv_2[26]), .B(n27839), .Y(n27838) );
  OAI211XL U31719 ( .A0(conv_2[26]), .A1(n27839), .B0(n27932), .C0(n27838), 
        .Y(n27840) );
  OAI211XL U31720 ( .A0(n30412), .A1(n27841), .B0(n33815), .C0(n27840), .Y(
        n15187) );
  AOI22XL U31721 ( .A0(n33620), .A1(n27843), .B0(n27842), .B1(n28673), .Y(
        n27845) );
  NAND2XL U31722 ( .A(n27847), .B(n27845), .Y(n27844) );
  OAI211XL U31723 ( .A0(n27847), .A1(n27845), .B0(n33778), .C0(n27844), .Y(
        n27846) );
  OAI211XL U31724 ( .A0(n30412), .A1(n27847), .B0(n35859), .C0(n27846), .Y(
        n15186) );
  NAND2XL U31725 ( .A(n27849), .B(n29046), .Y(n27853) );
  OAI21XL U31726 ( .A0(conv_2[198]), .A1(n27851), .B0(n27850), .Y(n27852) );
  NAND2XL U31727 ( .A(n27853), .B(n27852), .Y(n29041) );
  OAI21XL U31728 ( .A0(conv_2[199]), .A1(n29040), .B0(n29041), .Y(n27854) );
  NAND2XL U31729 ( .A(n35928), .B(n27854), .Y(n29941) );
  NAND2XL U31730 ( .A(conv_2[200]), .B(n29941), .Y(n35921) );
  NAND2XL U31731 ( .A(n29934), .B(conv_2[202]), .Y(n35927) );
  AOI21XL U31732 ( .A0(n29928), .A1(conv_2[204]), .B0(n29935), .Y(n29605) );
  NAND2XL U31733 ( .A(conv_2[205]), .B(n27856), .Y(n27855) );
  OAI211XL U31734 ( .A0(conv_2[205]), .A1(n27856), .B0(n32181), .C0(n27855), 
        .Y(n27857) );
  OAI211XL U31735 ( .A0(n35931), .A1(n27858), .B0(n34669), .C0(n27857), .Y(
        n15068) );
  NAND2XL U31736 ( .A(n29046), .B(n33509), .Y(n27866) );
  NAND2XL U31737 ( .A(n28068), .B(n33509), .Y(n27864) );
  OR2XL U31738 ( .A(n27859), .B(n18913), .Y(n27862) );
  NAND2XL U31739 ( .A(n27859), .B(n28126), .Y(n27861) );
  OAI22XL U31740 ( .A0(n27861), .A1(n27860), .B0(n27859), .B1(n28126), .Y(
        n30295) );
  NAND2XL U31741 ( .A(n30295), .B(conv_2[466]), .Y(n30294) );
  NAND2XL U31742 ( .A(n27862), .B(n30294), .Y(n30331) );
  AOI222XL U31743 ( .A0(n30332), .A1(conv_2[467]), .B0(n30332), .B1(n30331), 
        .C0(conv_2[467]), .C1(n30331), .Y(n27863) );
  NAND2XL U31744 ( .A(n27864), .B(n27863), .Y(n29560) );
  NAND2XL U31745 ( .A(n27866), .B(n27865), .Y(n28996) );
  NAND2XL U31746 ( .A(n27943), .B(n27867), .Y(n33891) );
  AOI21XL U31747 ( .A0(conv_2[470]), .A1(n33891), .B0(n34173), .Y(n27873) );
  NAND2XL U31748 ( .A(conv_2[471]), .B(n27869), .Y(n27868) );
  OAI211XL U31749 ( .A0(conv_2[471]), .A1(n27869), .B0(n33822), .C0(n27868), 
        .Y(n27870) );
  OAI211XL U31750 ( .A0(n34177), .A1(n27871), .B0(n34669), .C0(n27870), .Y(
        n14892) );
  NAND2XL U31751 ( .A(n27890), .B(n27885), .Y(n27879) );
  OAI2BB1XL U31752 ( .A0N(conv_2[472]), .A1N(n27886), .B0(n27943), .Y(n27880)
         );
  OAI2BB1XL U31753 ( .A0N(n34173), .A1N(n27879), .B0(n27880), .Y(n27876) );
  NAND2XL U31754 ( .A(n27878), .B(n27876), .Y(n27875) );
  OAI211XL U31755 ( .A0(n27878), .A1(n27876), .B0(n28751), .C0(n27875), .Y(
        n27877) );
  OAI211XL U31756 ( .A0(n34177), .A1(n27878), .B0(n34669), .C0(n27877), .Y(
        n14890) );
  AOI21XL U31757 ( .A0(conv_2[473]), .A1(n27880), .B0(n34173), .Y(n30900) );
  AOI21XL U31758 ( .A0(conv_2[475]), .A1(n34172), .B0(n34173), .Y(n27891) );
  INVXL U31759 ( .A(conv_2[475]), .Y(n34178) );
  NAND2XL U31760 ( .A(n34178), .B(n34171), .Y(n27892) );
  OAI21XL U31761 ( .A0(conv_2[476]), .A1(n27892), .B0(n34173), .Y(n27945) );
  OAI21XL U31762 ( .A0(n34173), .A1(n27944), .B0(n27945), .Y(n27883) );
  NAND2XL U31763 ( .A(n27946), .B(n27883), .Y(n27882) );
  OAI211XL U31764 ( .A0(n27946), .A1(n27883), .B0(n16656), .C0(n27882), .Y(
        n27884) );
  OAI211XL U31765 ( .A0(n34177), .A1(n27946), .B0(n34669), .C0(n27884), .Y(
        n14886) );
  OAI21XL U31766 ( .A0(n34173), .A1(n27886), .B0(n27885), .Y(n27888) );
  NAND2XL U31767 ( .A(n27890), .B(n27888), .Y(n27887) );
  OAI211XL U31768 ( .A0(n27890), .A1(n27888), .B0(n24499), .C0(n27887), .Y(
        n27889) );
  OAI211XL U31769 ( .A0(n34177), .A1(n27890), .B0(n34669), .C0(n27889), .Y(
        n14891) );
  AOI21XL U31770 ( .A0(n34173), .A1(n27892), .B0(n27891), .Y(n27894) );
  NAND2XL U31771 ( .A(conv_2[476]), .B(n27894), .Y(n27893) );
  OAI211XL U31772 ( .A0(conv_2[476]), .A1(n27894), .B0(n16656), .C0(n27893), 
        .Y(n27895) );
  OAI211XL U31773 ( .A0(n34177), .A1(n27896), .B0(n34669), .C0(n27895), .Y(
        n14887) );
  INVXL U31774 ( .A(conv_2[444]), .Y(n28795) );
  INVXL U31775 ( .A(conv_2[442]), .Y(n28941) );
  NAND2XL U31776 ( .A(n34224), .B(n28068), .Y(n27902) );
  NAND2XL U31777 ( .A(n34224), .B(n28128), .Y(n27900) );
  OAI21XL U31778 ( .A0(n27898), .A1(n18913), .B0(n27897), .Y(n30313) );
  OAI21XL U31779 ( .A0(conv_2[436]), .A1(n30312), .B0(n30313), .Y(n27899) );
  NAND2XL U31780 ( .A(n27900), .B(n27899), .Y(n30395) );
  OAI21XL U31781 ( .A0(conv_2[437]), .A1(n30394), .B0(n30395), .Y(n27901) );
  AND2XL U31782 ( .A(n27902), .B(n27901), .Y(n29554) );
  INVXL U31783 ( .A(conv_2[440]), .Y(n28947) );
  NAND2XL U31784 ( .A(conv_2[441]), .B(n36060), .Y(n28936) );
  NAND2XL U31785 ( .A(conv_2[443]), .B(n36066), .Y(n28791) );
  AOI2BB1XL U31786 ( .A0N(n36067), .A1N(n27921), .B0(n27922), .Y(n27907) );
  NAND2XL U31787 ( .A(conv_2[445]), .B(n27907), .Y(n27906) );
  OAI211XL U31788 ( .A0(conv_2[445]), .A1(n27907), .B0(n33778), .C0(n27906), 
        .Y(n27908) );
  OAI211XL U31789 ( .A0(n36070), .A1(n27909), .B0(n34669), .C0(n27908), .Y(
        n14908) );
  INVXL U31790 ( .A(conv_2[502]), .Y(n30910) );
  AOI21XL U31791 ( .A0(n36088), .A1(n30909), .B0(n30911), .Y(n27912) );
  NAND2XL U31792 ( .A(conv_2[502]), .B(n27912), .Y(n27911) );
  OAI211XL U31793 ( .A0(conv_2[502]), .A1(n27912), .B0(n34666), .C0(n27911), 
        .Y(n27913) );
  OAI211XL U31794 ( .A0(n36091), .A1(n30910), .B0(n34669), .C0(n27913), .Y(
        n14871) );
  AOI221XL U31795 ( .A0(n27915), .A1(n16656), .B0(n27914), .B1(n35336), .C0(
        n33615), .Y(n27920) );
  OAI211XL U31796 ( .A0(n33620), .A1(n27917), .B0(n34028), .C0(n27916), .Y(
        n27918) );
  OAI211XL U31797 ( .A0(n27920), .A1(n27919), .B0(n33815), .C0(n27918), .Y(
        n15188) );
  OAI2BB1XL U31798 ( .A0N(conv_2[445]), .A1N(n27921), .B0(n28937), .Y(n30961)
         );
  NAND4XL U31799 ( .A(conv_2[446]), .B(conv_2[447]), .C(n28937), .D(n30961), 
        .Y(n34731) );
  INVXL U31800 ( .A(conv_2[447]), .Y(n30966) );
  INVXL U31801 ( .A(conv_2[446]), .Y(n30870) );
  OAI21XL U31802 ( .A0(conv_2[445]), .A1(n27922), .B0(n36067), .Y(n30866) );
  NAND2XL U31803 ( .A(n30870), .B(n30866), .Y(n27923) );
  NAND3XL U31804 ( .A(n36067), .B(n30966), .C(n30962), .Y(n34730) );
  AOI22XL U31805 ( .A0(conv_2[448]), .A1(n34731), .B0(n34730), .B1(n34734), 
        .Y(n27925) );
  NAND2XL U31806 ( .A(conv_2[449]), .B(n27925), .Y(n27924) );
  OAI211XL U31807 ( .A0(conv_2[449]), .A1(n27925), .B0(n33788), .C0(n27924), 
        .Y(n27926) );
  OAI211XL U31808 ( .A0(n33442), .A1(n27927), .B0(n34669), .C0(n27926), .Y(
        n14904) );
  AOI22XL U31809 ( .A0(conv_2[13]), .A1(n27930), .B0(n27929), .B1(n27928), .Y(
        n27933) );
  NAND2XL U31810 ( .A(conv_2[14]), .B(n27933), .Y(n27931) );
  OAI211XL U31811 ( .A0(conv_2[14]), .A1(n27933), .B0(n27932), .C0(n27931), 
        .Y(n27934) );
  OAI211XL U31812 ( .A0(n33853), .A1(n27935), .B0(n35859), .C0(n27934), .Y(
        n15194) );
  AOI22XL U31813 ( .A0(conv_2[28]), .A1(n27938), .B0(n27937), .B1(n27936), .Y(
        n27940) );
  NAND2XL U31814 ( .A(conv_2[29]), .B(n27940), .Y(n27939) );
  OAI211XL U31815 ( .A0(conv_2[29]), .A1(n27940), .B0(n34666), .C0(n27939), 
        .Y(n27941) );
  OAI211XL U31816 ( .A0(n34676), .A1(n27942), .B0(n34669), .C0(n27941), .Y(
        n15184) );
  NAND3XL U31817 ( .A(n27944), .B(conv_2[477]), .C(n27943), .Y(n33275) );
  NAND3XL U31818 ( .A(n34173), .B(n27946), .C(n27945), .Y(n33274) );
  INVXL U31819 ( .A(conv_2[478]), .Y(n33278) );
  AOI22XL U31820 ( .A0(conv_2[478]), .A1(n33275), .B0(n33274), .B1(n33278), 
        .Y(n27948) );
  NAND2XL U31821 ( .A(conv_2[479]), .B(n27948), .Y(n27947) );
  OAI211XL U31822 ( .A0(conv_2[479]), .A1(n27948), .B0(n16656), .C0(n27947), 
        .Y(n27949) );
  OAI211XL U31823 ( .A0(n34520), .A1(n27950), .B0(n34669), .C0(n27949), .Y(
        n14884) );
  AOI22XL U31824 ( .A0(conv_2[43]), .A1(n27953), .B0(n27952), .B1(n27951), .Y(
        n27955) );
  NAND2XL U31825 ( .A(conv_2[44]), .B(n27955), .Y(n27954) );
  OAI211XL U31826 ( .A0(conv_2[44]), .A1(n27955), .B0(n16657), .C0(n27954), 
        .Y(n27956) );
  OAI211XL U31827 ( .A0(n33853), .A1(n27957), .B0(n34669), .C0(n27956), .Y(
        n15174) );
  AOI22XL U31828 ( .A0(conv_2[463]), .A1(n27960), .B0(n27959), .B1(n27958), 
        .Y(n27962) );
  NAND2XL U31829 ( .A(conv_2[464]), .B(n27962), .Y(n27961) );
  OAI211XL U31830 ( .A0(conv_2[464]), .A1(n27962), .B0(n32052), .C0(n27961), 
        .Y(n27963) );
  OAI211XL U31831 ( .A0(n34676), .A1(n27964), .B0(n34669), .C0(n27963), .Y(
        n14894) );
  INVXL U31832 ( .A(conv_1[283]), .Y(n29251) );
  ADDFX1 U31833 ( .A(conv_1[279]), .B(n29364), .CI(n27965), .CO(n29365), .S(
        n22288) );
  NAND4XL U31834 ( .A(conv_1[281]), .B(conv_1[282]), .C(n29339), .D(n35428), 
        .Y(n29253) );
  OAI21XL U31835 ( .A0(conv_1[280]), .A1(n29365), .B0(n29364), .Y(n35427) );
  NOR2BX1 U31836 ( .AN(n35427), .B(conv_1[281]), .Y(n35429) );
  INVXL U31837 ( .A(conv_1[282]), .Y(n29343) );
  NAND3XL U31838 ( .A(n35429), .B(n29364), .C(n29343), .Y(n29252) );
  NAND2XL U31839 ( .A(n29253), .B(n29252), .Y(n27968) );
  OAI21XL U31840 ( .A0(n16654), .A1(n27968), .B0(n35426), .Y(n27967) );
  NAND2XL U31841 ( .A(n27969), .B(n34281), .Y(n16180) );
  NAND2XL U31842 ( .A(conv_2[141]), .B(n30077), .Y(n35898) );
  NAND2XL U31843 ( .A(conv_2[143]), .B(n35906), .Y(n30088) );
  OAI2BB1XL U31844 ( .A0N(conv_2[145]), .A1N(n30095), .B0(n35899), .Y(n34357)
         );
  NAND4XL U31845 ( .A(conv_2[146]), .B(conv_2[147]), .C(n35899), .D(n34357), 
        .Y(n30235) );
  INVXL U31846 ( .A(conv_2[147]), .Y(n30086) );
  OAI21XL U31847 ( .A0(conv_2[145]), .A1(n30094), .B0(n35907), .Y(n34358) );
  NAND2XL U31848 ( .A(n34362), .B(n34358), .Y(n27973) );
  NAND3XL U31849 ( .A(n35907), .B(n30086), .C(n30082), .Y(n30234) );
  NAND2XL U31850 ( .A(n30235), .B(n30234), .Y(n27975) );
  OAI21XL U31851 ( .A0(n36009), .A1(n27975), .B0(n35902), .Y(n27974) );
  AOI32XL U31852 ( .A0(n36020), .A1(n30233), .A2(n27975), .B0(conv_2[148]), 
        .B1(n27974), .Y(n27976) );
  NAND2XL U31853 ( .A(n27976), .B(n35859), .Y(n15105) );
  AOI22XL U31854 ( .A0(n34808), .A1(n27978), .B0(n27977), .B1(n34810), .Y(
        N29234) );
  AOI22XL U31855 ( .A0(n34808), .A1(n27980), .B0(n27979), .B1(n34810), .Y(
        N29235) );
  AOI22XL U31856 ( .A0(conv_1[253]), .A1(n27983), .B0(n27982), .B1(n27981), 
        .Y(n27985) );
  NAND2XL U31857 ( .A(conv_1[254]), .B(n27985), .Y(n27984) );
  OAI211XL U31858 ( .A0(conv_1[254]), .A1(n27985), .B0(n33778), .C0(n27984), 
        .Y(n27986) );
  OAI211XL U31859 ( .A0(n33853), .A1(n27987), .B0(n16652), .C0(n27986), .Y(
        n16209) );
  INVXL U31860 ( .A(conv_3[390]), .Y(n27991) );
  AOI32XL U31861 ( .A0(n27988), .A1(n33703), .A2(n27990), .B0(n34389), .B1(
        n33703), .Y(n27989) );
  AOI32XL U31862 ( .A0(n34742), .A1(n27991), .A2(n27990), .B0(conv_3[390]), 
        .B1(n27989), .Y(n27992) );
  NAND2XL U31863 ( .A(n27992), .B(n34755), .Y(n15897) );
  ADDFXL U31864 ( .A(conv_2[351]), .B(n29526), .CI(n27993), .CO(n29523), .S(
        n23099) );
  INVXL U31865 ( .A(conv_2[352]), .Y(n29522) );
  NAND2XL U31866 ( .A(conv_2[353]), .B(n29525), .Y(n29480) );
  NAND2XL U31867 ( .A(n33925), .B(n29480), .Y(n27994) );
  INVXL U31868 ( .A(n27994), .Y(n27998) );
  NAND2XL U31869 ( .A(n29481), .B(n27995), .Y(n29479) );
  AOI32XL U31870 ( .A0(n27995), .A1(n36010), .A2(n27994), .B0(n16655), .B1(
        n36010), .Y(n27996) );
  AOI21XL U31871 ( .A0(conv_2[354]), .A1(n27996), .B0(n16651), .Y(n27997) );
  OAI31XL U31872 ( .A0(n27998), .A1(n16658), .A2(n29479), .B0(n27997), .Y(
        n14969) );
  AOI22XL U31873 ( .A0(conv_1[538]), .A1(n28001), .B0(n28000), .B1(n27999), 
        .Y(n28003) );
  NAND2XL U31874 ( .A(conv_1[539]), .B(n28003), .Y(n28002) );
  OAI211XL U31875 ( .A0(conv_1[539]), .A1(n28003), .B0(n24378), .C0(n28002), 
        .Y(n28004) );
  OAI211XL U31876 ( .A0(n33853), .A1(n28005), .B0(n34696), .C0(n28004), .Y(
        n15924) );
  NAND2XL U31877 ( .A(conv_2[275]), .B(n28009), .Y(n28008) );
  OAI211XL U31878 ( .A0(conv_2[275]), .A1(n28009), .B0(n16657), .C0(n28008), 
        .Y(n28010) );
  OAI211XL U31879 ( .A0(n30994), .A1(n28011), .B0(n33815), .C0(n28010), .Y(
        n15023) );
  NAND2XL U31880 ( .A(conv_2[384]), .B(n28015), .Y(n28014) );
  OAI211XL U31881 ( .A0(conv_2[384]), .A1(n28015), .B0(n32611), .C0(n28014), 
        .Y(n28016) );
  OAI211XL U31882 ( .A0(n36028), .A1(n28017), .B0(n34669), .C0(n28016), .Y(
        n14949) );
  INVXL U31883 ( .A(conv_2[387]), .Y(n28022) );
  ADDFX1 U31884 ( .A(conv_2[385]), .B(n34529), .CI(n28018), .CO(n34528), .S(
        n23080) );
  INVXL U31885 ( .A(conv_2[386]), .Y(n34533) );
  OAI33XL U31886 ( .A0(conv_2[386]), .A1(n34528), .A2(n36025), .B0(n34533), 
        .B1(n34537), .B2(n34529), .Y(n28020) );
  NAND2XL U31887 ( .A(conv_2[387]), .B(n28020), .Y(n28019) );
  OAI211XL U31888 ( .A0(conv_2[387]), .A1(n28020), .B0(n16657), .C0(n28019), 
        .Y(n28021) );
  OAI211XL U31889 ( .A0(n36028), .A1(n28022), .B0(n33815), .C0(n28021), .Y(
        n14946) );
  INVXL U31890 ( .A(conv_2[279]), .Y(n28040) );
  OAI2BB1XL U31891 ( .A0N(conv_2[277]), .A1N(n28767), .B0(n28883), .Y(n28032)
         );
  NAND2XL U31892 ( .A(conv_2[278]), .B(n28032), .Y(n28039) );
  INVXL U31893 ( .A(conv_2[277]), .Y(n28771) );
  NAND2XL U31894 ( .A(n35950), .B(n28025), .Y(n28766) );
  NAND2XL U31895 ( .A(n28771), .B(n28766), .Y(n28033) );
  AOI21XL U31896 ( .A0(n28883), .A1(n28039), .B0(n28038), .Y(n28027) );
  NAND2XL U31897 ( .A(conv_2[279]), .B(n28027), .Y(n28026) );
  OAI211XL U31898 ( .A0(conv_2[279]), .A1(n28027), .B0(n33778), .C0(n28026), 
        .Y(n28028) );
  OAI211XL U31899 ( .A0(n30994), .A1(n28040), .B0(n34669), .C0(n28028), .Y(
        n15019) );
  INVXL U31900 ( .A(conv_2[388]), .Y(n28154) );
  NAND4XL U31901 ( .A(conv_2[386]), .B(conv_2[387]), .C(n34528), .D(n36025), 
        .Y(n28156) );
  NAND2XL U31902 ( .A(n28156), .B(n28155), .Y(n28030) );
  NAND2XL U31903 ( .A(conv_2[388]), .B(n28030), .Y(n28029) );
  OAI211XL U31904 ( .A0(conv_2[388]), .A1(n28030), .B0(n33788), .C0(n28029), 
        .Y(n28031) );
  OAI211XL U31905 ( .A0(n36028), .A1(n28154), .B0(n35859), .C0(n28031), .Y(
        n14945) );
  INVXL U31906 ( .A(conv_2[278]), .Y(n28037) );
  OAI2BB1XL U31907 ( .A0N(n35950), .A1N(n28033), .B0(n28032), .Y(n28035) );
  NAND2XL U31908 ( .A(n28037), .B(n28035), .Y(n28034) );
  OAI211XL U31909 ( .A0(n28037), .A1(n28035), .B0(n33788), .C0(n28034), .Y(
        n28036) );
  OAI211XL U31910 ( .A0(n30994), .A1(n28037), .B0(n34735), .C0(n28036), .Y(
        n15020) );
  INVXL U31911 ( .A(conv_2[281]), .Y(n28885) );
  AOI2BB1XL U31912 ( .A0N(conv_2[279]), .A1N(n28038), .B0(n28883), .Y(n35948)
         );
  OAI21XL U31913 ( .A0(conv_2[280]), .A1(n35948), .B0(n35950), .Y(n28884) );
  OAI2BB1XL U31914 ( .A0N(conv_2[280]), .A1N(n35949), .B0(n28883), .Y(n30985)
         );
  NAND2XL U31915 ( .A(n28884), .B(n30985), .Y(n28042) );
  NAND2XL U31916 ( .A(n28885), .B(n28042), .Y(n28041) );
  OAI211XL U31917 ( .A0(n28885), .A1(n28042), .B0(n32656), .C0(n28041), .Y(
        n28043) );
  OAI211XL U31918 ( .A0(n30994), .A1(n28885), .B0(n34735), .C0(n28043), .Y(
        n15017) );
  INVXL U31919 ( .A(conv_2[323]), .Y(n28049) );
  AOI2BB1XL U31920 ( .A0N(conv_2[322]), .A1N(n35983), .B0(n33079), .Y(n28044)
         );
  AOI2BB1XL U31921 ( .A0N(n35982), .A1N(n28045), .B0(n28044), .Y(n28047) );
  NAND2XL U31922 ( .A(conv_2[323]), .B(n28047), .Y(n28046) );
  OAI211XL U31923 ( .A0(conv_2[323]), .A1(n28047), .B0(n30090), .C0(n28046), 
        .Y(n28048) );
  OAI211XL U31924 ( .A0(n35986), .A1(n28049), .B0(n34735), .C0(n28048), .Y(
        n14990) );
  INVXL U31925 ( .A(conv_2[320]), .Y(n28055) );
  NAND2XL U31926 ( .A(conv_2[320]), .B(n28053), .Y(n28052) );
  OAI211XL U31927 ( .A0(conv_2[320]), .A1(n28053), .B0(n33982), .C0(n28052), 
        .Y(n28054) );
  OAI211XL U31928 ( .A0(n35986), .A1(n28055), .B0(n35859), .C0(n28054), .Y(
        n14993) );
  INVXL U31929 ( .A(conv_2[325]), .Y(n28062) );
  NAND2XL U31930 ( .A(conv_2[325]), .B(n28060), .Y(n28059) );
  OAI211XL U31931 ( .A0(conv_2[325]), .A1(n28060), .B0(n30090), .C0(n28059), 
        .Y(n28061) );
  OAI211XL U31932 ( .A0(n35986), .A1(n28062), .B0(n34735), .C0(n28061), .Y(
        n14988) );
  INVXL U31933 ( .A(conv_2[326]), .Y(n33081) );
  OAI21XL U31934 ( .A0(conv_2[325]), .A1(n28063), .B0(n35982), .Y(n33080) );
  NAND2XL U31935 ( .A(n33080), .B(n33933), .Y(n28066) );
  NAND2XL U31936 ( .A(n33081), .B(n28066), .Y(n28065) );
  OAI211XL U31937 ( .A0(n33081), .A1(n28066), .B0(n33788), .C0(n28065), .Y(
        n28067) );
  OAI211XL U31938 ( .A0(n35986), .A1(n33081), .B0(n34669), .C0(n28067), .Y(
        n14987) );
  INVXL U31939 ( .A(conv_2[412]), .Y(n28080) );
  NAND2XL U31940 ( .A(n29046), .B(n34229), .Y(n28075) );
  NAND2XL U31941 ( .A(n28068), .B(n34229), .Y(n28073) );
  OR2XL U31942 ( .A(n28069), .B(n18913), .Y(n29794) );
  OAI21XL U31943 ( .A0(n18913), .A1(n28070), .B0(n28069), .Y(n29793) );
  NAND2XL U31944 ( .A(conv_2[406]), .B(n29793), .Y(n28071) );
  NAND2XL U31945 ( .A(n29794), .B(n28071), .Y(n29965) );
  AOI222XL U31946 ( .A0(n29966), .A1(conv_2[407]), .B0(n29966), .B1(n29965), 
        .C0(conv_2[407]), .C1(n29965), .Y(n28072) );
  NAND2XL U31947 ( .A(n28073), .B(n28072), .Y(n29421) );
  NAND2XL U31948 ( .A(n28075), .B(n28074), .Y(n28859) );
  NAND2XL U31949 ( .A(n33321), .B(n28076), .Y(n33379) );
  NAND2XL U31950 ( .A(conv_2[410]), .B(n33379), .Y(n29487) );
  AOI2BB1XL U31951 ( .A0N(n36045), .A1N(n28081), .B0(n28082), .Y(n28078) );
  NAND2XL U31952 ( .A(conv_2[412]), .B(n28078), .Y(n28077) );
  OAI211XL U31953 ( .A0(conv_2[412]), .A1(n28078), .B0(n33788), .C0(n28077), 
        .Y(n28079) );
  OAI211XL U31954 ( .A0(n36047), .A1(n28080), .B0(n33815), .C0(n28079), .Y(
        n14931) );
  NAND2XL U31955 ( .A(n28081), .B(conv_2[412]), .Y(n30885) );
  AOI21XL U31956 ( .A0(n33321), .A1(n30885), .B0(n30883), .Y(n28084) );
  NAND2XL U31957 ( .A(conv_2[413]), .B(n28084), .Y(n28083) );
  OAI211XL U31958 ( .A0(conv_2[413]), .A1(n28084), .B0(n33788), .C0(n28083), 
        .Y(n28085) );
  OAI211XL U31959 ( .A0(n36047), .A1(n30884), .B0(n34669), .C0(n28085), .Y(
        n14930) );
  INVXL U31960 ( .A(conv_2[292]), .Y(n28095) );
  INVXL U31961 ( .A(n28088), .Y(n28089) );
  INVXL U31962 ( .A(conv_2[290]), .Y(n30892) );
  AOI21XL U31963 ( .A0(n35956), .A1(conv_2[291]), .B0(n35957), .Y(n30916) );
  NAND2XL U31964 ( .A(conv_2[292]), .B(n28093), .Y(n28092) );
  OAI211XL U31965 ( .A0(conv_2[292]), .A1(n28093), .B0(n24378), .C0(n28092), 
        .Y(n28094) );
  OAI211XL U31966 ( .A0(n35963), .A1(n28095), .B0(n34669), .C0(n28094), .Y(
        n15011) );
  INVXL U31967 ( .A(conv_2[335]), .Y(n28101) );
  NOR2BXL U31968 ( .AN(n28097), .B(n28096), .Y(n28099) );
  NAND2XL U31969 ( .A(conv_2[335]), .B(n28099), .Y(n28098) );
  OAI211XL U31970 ( .A0(conv_2[335]), .A1(n28099), .B0(n32611), .C0(n28098), 
        .Y(n28100) );
  OAI211XL U31971 ( .A0(n36003), .A1(n28101), .B0(n34735), .C0(n28100), .Y(
        n14983) );
  INVXL U31972 ( .A(conv_2[338]), .Y(n28107) );
  ADDFXL U31973 ( .A(conv_2[337]), .B(n35995), .CI(n28102), .CO(n35996), .S(
        n23087) );
  AOI21XL U31974 ( .A0(n35996), .A1(n35995), .B0(n28103), .Y(n28105) );
  NAND2XL U31975 ( .A(conv_2[338]), .B(n28105), .Y(n28104) );
  OAI211XL U31976 ( .A0(conv_2[338]), .A1(n28105), .B0(n33982), .C0(n28104), 
        .Y(n28106) );
  OAI211XL U31977 ( .A0(n36003), .A1(n28107), .B0(n34735), .C0(n28106), .Y(
        n14980) );
  NAND2XL U31978 ( .A(conv_2[396]), .B(n28111), .Y(n28110) );
  OAI211XL U31979 ( .A0(conv_2[396]), .A1(n28111), .B0(n33788), .C0(n28110), 
        .Y(n28112) );
  OAI211XL U31980 ( .A0(n36031), .A1(n28113), .B0(n35859), .C0(n28112), .Y(
        n14942) );
  NAND2XL U31981 ( .A(conv_2[395]), .B(n28117), .Y(n28116) );
  OAI211XL U31982 ( .A0(conv_2[395]), .A1(n28117), .B0(n24378), .C0(n28116), 
        .Y(n28118) );
  OAI211XL U31983 ( .A0(n36031), .A1(n28119), .B0(n33815), .C0(n28118), .Y(
        n14943) );
  INVXL U31984 ( .A(conv_2[357]), .Y(n29461) );
  OAI2BB1XL U31985 ( .A0N(conv_2[355]), .A1N(n28120), .B0(n33925), .Y(n36012)
         );
  OAI21XL U31986 ( .A0(conv_2[355]), .A1(n29479), .B0(n29526), .Y(n36011) );
  AOI32XL U31987 ( .A0(conv_2[356]), .A1(n33925), .A2(n36012), .B0(n29526), 
        .B1(n36013), .Y(n28122) );
  NAND2XL U31988 ( .A(n29461), .B(n28122), .Y(n28121) );
  OAI211XL U31989 ( .A0(n29461), .A1(n28122), .B0(n32181), .C0(n28121), .Y(
        n28123) );
  OAI211XL U31990 ( .A0(n36010), .A1(n29461), .B0(n34735), .C0(n28123), .Y(
        n14966) );
  INVXL U31991 ( .A(conv_2[425]), .Y(n28891) );
  INVXL U31992 ( .A(conv_2[421]), .Y(n29820) );
  NAND2XL U31993 ( .A(n28124), .B(conv_2[420]), .Y(n28125) );
  OAI2BB1XL U31994 ( .A0N(n28125), .A1N(n18913), .B0(n34768), .Y(n29815) );
  NAND2XL U31995 ( .A(n34488), .B(n28126), .Y(n29816) );
  NAND2XL U31996 ( .A(n35853), .B(n28129), .Y(n28127) );
  OAI31XL U31997 ( .A0(n35853), .A1(n35499), .A2(n28129), .B0(n28127), .Y(
        n30011) );
  NAND2XL U31998 ( .A(n28129), .B(n28128), .Y(n28130) );
  OAI2BB1XL U31999 ( .A0N(conv_2[422]), .A1N(n30011), .B0(n28130), .Y(n32870)
         );
  NAND2XL U32000 ( .A(conv_2[425]), .B(n28135), .Y(n28134) );
  OAI211XL U32001 ( .A0(conv_2[425]), .A1(n28135), .B0(n32052), .C0(n28134), 
        .Y(n28136) );
  OAI211XL U32002 ( .A0(n36053), .A1(n28891), .B0(n34735), .C0(n28136), .Y(
        n14923) );
  OAI2BB1XL U32003 ( .A0N(n28138), .A1N(conv_2[264]), .B0(n28161), .Y(n28184)
         );
  OAI31XL U32004 ( .A0(conv_2[263]), .A1(conv_2[264]), .A2(n28190), .B0(n28191), .Y(n28183) );
  NAND2XL U32005 ( .A(n28188), .B(n28183), .Y(n28167) );
  NAND2XL U32006 ( .A(n28184), .B(n28167), .Y(n28140) );
  NAND2XL U32007 ( .A(n28161), .B(n28140), .Y(n28166) );
  AND2XL U32008 ( .A(n28140), .B(n28171), .Y(n28139) );
  AOI32XL U32009 ( .A0(conv_2[266]), .A1(n28166), .A2(n28161), .B0(n28139), 
        .B1(n28166), .Y(n28174) );
  NAND2XL U32010 ( .A(n28172), .B(n28161), .Y(n28197) );
  NAND4XL U32011 ( .A(n28171), .B(n28140), .C(n28176), .D(n28191), .Y(n28196)
         );
  AOI22XL U32012 ( .A0(conv_2[268]), .A1(n28197), .B0(n28196), .B1(n28201), 
        .Y(n28142) );
  NAND2XL U32013 ( .A(conv_2[269]), .B(n28142), .Y(n28141) );
  OAI211XL U32014 ( .A0(conv_2[269]), .A1(n28142), .B0(n35336), .C0(n28141), 
        .Y(n28143) );
  OAI211XL U32015 ( .A0(n34676), .A1(n28144), .B0(n34735), .C0(n28143), .Y(
        n15024) );
  NAND2XL U32016 ( .A(n29046), .B(n33535), .Y(n28148) );
  NAND2XL U32017 ( .A(n28148), .B(n28147), .Y(n28978) );
  NAND2XL U32018 ( .A(n29455), .B(n28149), .Y(n28259) );
  NAND2XL U32019 ( .A(conv_2[245]), .B(n28259), .Y(n29144) );
  NAND2XL U32020 ( .A(conv_2[247]), .B(n29168), .Y(n29150) );
  INVXL U32021 ( .A(n29455), .Y(n35942) );
  AOI21XL U32022 ( .A0(conv_2[249]), .A1(n33683), .B0(n35942), .Y(n33199) );
  OAI2BB1XL U32023 ( .A0N(conv_2[251]), .A1N(n35941), .B0(n29455), .Y(n29454)
         );
  NAND3XL U32024 ( .A(conv_2[252]), .B(n29455), .C(n29454), .Y(n34145) );
  NAND3XL U32025 ( .A(n35942), .B(n29456), .C(n29460), .Y(n34144) );
  AOI22XL U32026 ( .A0(conv_2[253]), .A1(n34145), .B0(n34144), .B1(n34148), 
        .Y(n28151) );
  NAND2XL U32027 ( .A(conv_2[254]), .B(n28151), .Y(n28150) );
  OAI211XL U32028 ( .A0(conv_2[254]), .A1(n28151), .B0(n35336), .C0(n28150), 
        .Y(n28152) );
  OAI211XL U32029 ( .A0(n34520), .A1(n28153), .B0(n35859), .C0(n28152), .Y(
        n15034) );
  NAND2XL U32030 ( .A(conv_2[389]), .B(n28158), .Y(n28157) );
  OAI211XL U32031 ( .A0(conv_2[389]), .A1(n28158), .B0(n27932), .C0(n28157), 
        .Y(n28159) );
  OAI33XL U32032 ( .A0(conv_2[263]), .A1(n28161), .A2(n28190), .B0(n28195), 
        .B1(n28189), .B2(n28191), .Y(n28163) );
  NAND2XL U32033 ( .A(conv_2[264]), .B(n28163), .Y(n28162) );
  OAI211XL U32034 ( .A0(conv_2[264]), .A1(n28163), .B0(n33778), .C0(n28162), 
        .Y(n28164) );
  OAI211XL U32035 ( .A0(n34601), .A1(n28165), .B0(n33815), .C0(n28164), .Y(
        n15029) );
  OAI2BB1XL U32036 ( .A0N(n28191), .A1N(n28167), .B0(n28166), .Y(n28169) );
  NAND2XL U32037 ( .A(n28171), .B(n28169), .Y(n28168) );
  OAI211XL U32038 ( .A0(n28171), .A1(n28169), .B0(n28751), .C0(n28168), .Y(
        n28170) );
  OAI211XL U32039 ( .A0(n34601), .A1(n28171), .B0(n34669), .C0(n28170), .Y(
        n15027) );
  OAI2BB1XL U32040 ( .A0N(n28176), .A1N(n28174), .B0(n28173), .Y(n28175) );
  OAI211XL U32041 ( .A0(n34601), .A1(n28176), .B0(n34735), .C0(n28175), .Y(
        n15026) );
  NAND2XL U32042 ( .A(conv_2[260]), .B(n28180), .Y(n28179) );
  OAI211XL U32043 ( .A0(conv_2[260]), .A1(n28180), .B0(n16657), .C0(n28179), 
        .Y(n28181) );
  OAI211XL U32044 ( .A0(n34601), .A1(n28182), .B0(n34735), .C0(n28181), .Y(
        n15033) );
  NAND2XL U32045 ( .A(n28184), .B(n28183), .Y(n28186) );
  NAND2XL U32046 ( .A(n28188), .B(n28186), .Y(n28185) );
  OAI211XL U32047 ( .A0(n28188), .A1(n28186), .B0(n28751), .C0(n28185), .Y(
        n28187) );
  OAI211XL U32048 ( .A0(n34601), .A1(n28188), .B0(n35859), .C0(n28187), .Y(
        n15028) );
  AOI21XL U32049 ( .A0(n28191), .A1(n28190), .B0(n28189), .Y(n28193) );
  NAND2XL U32050 ( .A(conv_2[263]), .B(n28193), .Y(n28192) );
  OAI211XL U32051 ( .A0(conv_2[263]), .A1(n28193), .B0(n34028), .C0(n28192), 
        .Y(n28194) );
  OAI211XL U32052 ( .A0(n34601), .A1(n28195), .B0(n33815), .C0(n28194), .Y(
        n15030) );
  NAND2XL U32053 ( .A(n28197), .B(n28196), .Y(n28199) );
  NAND2XL U32054 ( .A(conv_2[268]), .B(n28199), .Y(n28198) );
  OAI211XL U32055 ( .A0(conv_2[268]), .A1(n28199), .B0(n35336), .C0(n28198), 
        .Y(n28200) );
  OAI211XL U32056 ( .A0(n34601), .A1(n28201), .B0(n34669), .C0(n28200), .Y(
        n15025) );
  NAND4XL U32057 ( .A(conv_2[521]), .B(conv_2[522]), .C(n28706), .D(n31008), 
        .Y(n29439) );
  NAND3XL U32058 ( .A(n33580), .B(n28203), .C(n28202), .Y(n29438) );
  NAND2XL U32059 ( .A(n29439), .B(n29438), .Y(n28205) );
  NAND2XL U32060 ( .A(conv_2[523]), .B(n28205), .Y(n28204) );
  OAI211XL U32061 ( .A0(conv_2[523]), .A1(n28205), .B0(n33982), .C0(n28204), 
        .Y(n28206) );
  OAI211XL U32062 ( .A0(n31013), .A1(n29437), .B0(n34669), .C0(n28206), .Y(
        n14855) );
  OAI2BB1XL U32063 ( .A0N(n28211), .A1N(n28210), .B0(n28209), .Y(n33336) );
  AOI22XL U32064 ( .A0(affine_2[46]), .A1(n33367), .B0(n16674), .B1(n28214), 
        .Y(n28215) );
  NAND2XL U32065 ( .A(n28215), .B(n33340), .Y(n16547) );
  AOI22XL U32066 ( .A0(n36120), .A1(n28217), .B0(n28216), .B1(n28249), .Y(
        n14675) );
  INVXL U32067 ( .A(filter_1[49]), .Y(n28219) );
  INVXL U32068 ( .A(filter_1[43]), .Y(n28224) );
  AOI22XL U32069 ( .A0(n36120), .A1(n28219), .B0(n28224), .B1(n28249), .Y(
        n14707) );
  INVXL U32070 ( .A(filter_1[29]), .Y(n28226) );
  AOI22XL U32071 ( .A0(n36120), .A1(n28226), .B0(n28218), .B1(n28249), .Y(
        n14667) );
  INVXL U32072 ( .A(filter_1[52]), .Y(n28222) );
  AOI22XL U32073 ( .A0(n36120), .A1(n36148), .B0(n28222), .B1(n28249), .Y(
        n14681) );
  AOI22XL U32074 ( .A0(n36120), .A1(n36139), .B0(n28219), .B1(n28249), .Y(
        n14708) );
  INVXL U32075 ( .A(filter_1[24]), .Y(n28239) );
  AOI22XL U32076 ( .A0(n36120), .A1(n28220), .B0(n28239), .B1(n28249), .Y(
        n14713) );
  AOI22XL U32077 ( .A0(n36120), .A1(n28222), .B0(n28221), .B1(n28249), .Y(
        n14680) );
  INVXL U32078 ( .A(filter_1[12]), .Y(n28235) );
  INVXL U32079 ( .A(filter_1[6]), .Y(n36115) );
  AOI22XL U32080 ( .A0(n36120), .A1(n28235), .B0(n36115), .B1(n28249), .Y(
        n14710) );
  INVXL U32081 ( .A(filter_1[15]), .Y(n28225) );
  INVXL U32082 ( .A(filter_1[9]), .Y(n36118) );
  AOI22XL U32083 ( .A0(n36120), .A1(n28225), .B0(n36118), .B1(n28249), .Y(
        n14683) );
  INVXL U32084 ( .A(filter_1[42]), .Y(n28229) );
  AOI22XL U32085 ( .A0(n36120), .A1(n28223), .B0(n28229), .B1(n28249), .Y(
        n14716) );
  INVXL U32086 ( .A(filter_1[37]), .Y(n28251) );
  AOI22XL U32087 ( .A0(n36120), .A1(n28224), .B0(n28251), .B1(n28249), .Y(
        n14706) );
  INVXL U32088 ( .A(filter_1[21]), .Y(n28246) );
  AOI22XL U32089 ( .A0(n36120), .A1(n28246), .B0(n28225), .B1(n28249), .Y(
        n14684) );
  AOI22XL U32090 ( .A0(n36120), .A1(n28227), .B0(n28226), .B1(n28249), .Y(
        n14668) );
  AOI22XL U32091 ( .A0(n36120), .A1(n28229), .B0(n28228), .B1(n28249), .Y(
        n14715) );
  INVXL U32092 ( .A(filter_1[33]), .Y(n28232) );
  INVXL U32093 ( .A(filter_1[27]), .Y(n28247) );
  AOI22XL U32094 ( .A0(n36120), .A1(n28232), .B0(n28247), .B1(n28249), .Y(
        n14686) );
  AOI22XL U32095 ( .A0(n36120), .A1(n28231), .B0(n28230), .B1(n28249), .Y(
        n14677) );
  AOI22XL U32096 ( .A0(n36120), .A1(n28233), .B0(n28232), .B1(n28249), .Y(
        n14687) );
  INVXL U32097 ( .A(filter_1[8]), .Y(n36117) );
  AOI22XL U32098 ( .A0(n36120), .A1(n28234), .B0(n36117), .B1(n28249), .Y(
        n14692) );
  INVXL U32099 ( .A(filter_1[18]), .Y(n28238) );
  AOI22XL U32100 ( .A0(n36120), .A1(n28238), .B0(n28235), .B1(n28249), .Y(
        n14711) );
  INVXL U32101 ( .A(filter_1[26]), .Y(n28237) );
  AOI22XL U32102 ( .A0(n36120), .A1(n28237), .B0(n28236), .B1(n28249), .Y(
        n14694) );
  INVXL U32103 ( .A(filter_1[32]), .Y(n28240) );
  AOI22XL U32104 ( .A0(n36120), .A1(n28240), .B0(n28237), .B1(n28249), .Y(
        n14695) );
  AOI22XL U32105 ( .A0(n36120), .A1(n28239), .B0(n28238), .B1(n28249), .Y(
        n14712) );
  INVXL U32106 ( .A(filter_1[38]), .Y(n28241) );
  AOI22XL U32107 ( .A0(n36120), .A1(n28241), .B0(n28240), .B1(n28249), .Y(
        n14696) );
  INVXL U32108 ( .A(filter_1[44]), .Y(n28242) );
  AOI22XL U32109 ( .A0(n36120), .A1(n28242), .B0(n28241), .B1(n28249), .Y(
        n14697) );
  INVXL U32110 ( .A(filter_1[50]), .Y(n28243) );
  AOI22XL U32111 ( .A0(n36120), .A1(n28243), .B0(n28242), .B1(n28249), .Y(
        n14698) );
  AOI22XL U32112 ( .A0(n36120), .A1(n36142), .B0(n28243), .B1(n28249), .Y(
        n14699) );
  INVXL U32113 ( .A(filter_1[13]), .Y(n28244) );
  INVXL U32114 ( .A(filter_1[7]), .Y(n36116) );
  AOI22XL U32115 ( .A0(n36120), .A1(n28244), .B0(n36116), .B1(n28249), .Y(
        n14701) );
  INVXL U32116 ( .A(filter_1[19]), .Y(n28245) );
  AOI22XL U32117 ( .A0(n36120), .A1(n28245), .B0(n28244), .B1(n28249), .Y(
        n14702) );
  INVXL U32118 ( .A(filter_1[25]), .Y(n28248) );
  AOI22XL U32119 ( .A0(n36120), .A1(n28248), .B0(n28245), .B1(n28249), .Y(
        n14703) );
  AOI22XL U32120 ( .A0(n36120), .A1(n28247), .B0(n28246), .B1(n28249), .Y(
        n14685) );
  INVXL U32121 ( .A(filter_1[31]), .Y(n28250) );
  AOI22XL U32122 ( .A0(n36120), .A1(n28250), .B0(n28248), .B1(n28249), .Y(
        n14704) );
  AOI22XL U32123 ( .A0(n36120), .A1(n28251), .B0(n28250), .B1(n28249), .Y(
        n14705) );
  NAND3XL U32124 ( .A(n28252), .B(conv_2[537]), .C(n29095), .Y(n30423) );
  NAND3XL U32125 ( .A(n28254), .B(n33629), .C(n28253), .Y(n30422) );
  NAND2XL U32126 ( .A(n30423), .B(n30422), .Y(n28256) );
  NAND2XL U32127 ( .A(conv_2[538]), .B(n28256), .Y(n28255) );
  OAI211XL U32128 ( .A0(conv_2[538]), .A1(n28256), .B0(n32052), .C0(n28255), 
        .Y(n28257) );
  OAI211XL U32129 ( .A0(n34496), .A1(n30421), .B0(n34735), .C0(n28257), .Y(
        n14845) );
  NOR2BXL U32130 ( .AN(n28259), .B(n28258), .Y(n28261) );
  NAND2XL U32131 ( .A(conv_2[245]), .B(n28261), .Y(n28260) );
  OAI211XL U32132 ( .A0(conv_2[245]), .A1(n28261), .B0(n32052), .C0(n28260), 
        .Y(n28262) );
  OAI211XL U32133 ( .A0(n35945), .A1(n28263), .B0(n34735), .C0(n28262), .Y(
        n15043) );
  OAI2BB2X1 U32134 ( .B0(n35170), .B1(n28349), .A0N(n35167), .A1N(n34963), .Y(
        n28269) );
  AOI22XL U32135 ( .A0(n16665), .A1(n28264), .B0(n35169), .B1(n28372), .Y(
        n28267) );
  AOI22XL U32136 ( .A0(n28324), .A1(n35168), .B0(n28559), .B1(n28265), .Y(
        n28266) );
  OAI211XL U32137 ( .A0(n35171), .A1(n18196), .B0(n28267), .C0(n28266), .Y(
        n28268) );
  INVXL U32138 ( .A(pool[108]), .Y(n35009) );
  OAI21XL U32139 ( .A0(n35126), .A1(n26621), .B0(n28270), .Y(n28272) );
  OAI22XL U32140 ( .A0(n35136), .A1(n34989), .B0(n16701), .B1(n35134), .Y(
        n28271) );
  OAI2BB1XL U32141 ( .A0N(n16670), .A1N(n35140), .B0(n28275), .Y(n28284) );
  OAI2BB2XL U32142 ( .B0(n35141), .B1(n28575), .A0N(n35148), .A1N(n28324), .Y(
        n28283) );
  OAI22XL U32143 ( .A0(n35142), .A1(n28277), .B0(n28276), .B1(n28349), .Y(
        n28282) );
  AOI222XL U32144 ( .A0(n28280), .A1(n28291), .B0(n28279), .B1(n28290), .C0(
        n28278), .C1(n28289), .Y(n35145) );
  OAI22XL U32145 ( .A0(n35145), .A1(n28467), .B0(n16701), .B1(n35144), .Y(
        n28281) );
  AOI2BB2XL U32146 ( .B0(n16665), .B1(n35235), .A0N(n26621), .A1N(n35240), .Y(
        n28287) );
  INVXL U32147 ( .A(n28285), .Y(n35233) );
  OAI211XL U32148 ( .A0(n34982), .A1(n28304), .B0(n28287), .C0(n28286), .Y(
        n28296) );
  INVXL U32149 ( .A(n28288), .Y(n34985) );
  AOI222XL U32150 ( .A0(n34986), .A1(n28291), .B0(n34985), .B1(n28290), .C0(
        n35230), .C1(n28289), .Y(n35243) );
  AOI22XL U32151 ( .A0(n36245), .A1(n28294), .B0(n28293), .B1(n28292), .Y(
        n35242) );
  OAI22XL U32152 ( .A0(n35243), .A1(n28467), .B0(n16701), .B1(n35242), .Y(
        n28295) );
  AOI22XL U32153 ( .A0(n16665), .A1(n35154), .B0(n28366), .B1(n35152), .Y(
        n28300) );
  OAI22XL U32154 ( .A0(n35160), .A1(n34989), .B0(n16701), .B1(n35158), .Y(
        n28297) );
  AOI222XL U32155 ( .A0(n35003), .A1(n35005), .B0(n35003), .B1(n35004), .C0(
        n35005), .C1(n35004), .Y(n28302) );
  AOI222XL U32156 ( .A0(n35007), .A1(pool[107]), .B0(n35007), .B1(n28302), 
        .C0(pool[107]), .C1(n28302), .Y(n28303) );
  OAI22XL U32157 ( .A0(n24828), .A1(n28304), .B0(n35103), .B1(n28349), .Y(
        n28306) );
  OAI22XL U32158 ( .A0(n35109), .A1(n34989), .B0(n16701), .B1(n35108), .Y(
        n28305) );
  NAND2XL U32159 ( .A(n16670), .B(n35102), .Y(n28307) );
  OAI211XL U32160 ( .A0(n35107), .A1(n26621), .B0(n28308), .C0(n28307), .Y(
        n28338) );
  AOI22XL U32161 ( .A0(n28366), .A1(n35052), .B0(n16663), .B1(n35044), .Y(
        n28314) );
  OAI22XL U32162 ( .A0(n28310), .A1(n28575), .B0(n28309), .B1(n28333), .Y(
        n28312) );
  OAI22XL U32163 ( .A0(n35042), .A1(n16672), .B0(n35041), .B1(n28553), .Y(
        n28311) );
  AOI211XL U32164 ( .A0(n34961), .A1(n35043), .B0(n28312), .C0(n28311), .Y(
        n28313) );
  OAI211XL U32165 ( .A0(n26575), .A1(n35049), .B0(n28314), .C0(n28313), .Y(
        n28328) );
  AOI22XL U32166 ( .A0(n28366), .A1(n35092), .B0(n18463), .B1(n35094), .Y(
        n28320) );
  OAI22XL U32167 ( .A0(n28316), .A1(n28575), .B0(n28315), .B1(n28349), .Y(
        n28318) );
  OAI22XL U32168 ( .A0(n35090), .A1(n28333), .B0(n35089), .B1(n18196), .Y(
        n28317) );
  AOI211XL U32169 ( .A0(n16665), .A1(n35091), .B0(n28318), .C0(n28317), .Y(
        n28319) );
  OAI211XL U32170 ( .A0(n26575), .A1(n35097), .B0(n28320), .C0(n28319), .Y(
        n28327) );
  AOI22XL U32171 ( .A0(n28414), .A1(n35069), .B0(n34961), .B1(n35066), .Y(
        n28326) );
  OAI22XL U32172 ( .A0(n35068), .A1(n16672), .B0(n35067), .B1(n28553), .Y(
        n28323) );
  OAI22XL U32173 ( .A0(n35070), .A1(n28333), .B0(n35065), .B1(n28349), .Y(
        n28322) );
  AOI211XL U32174 ( .A0(n28324), .A1(n35073), .B0(n28323), .C0(n28322), .Y(
        n28325) );
  OAI211XL U32175 ( .A0(n26575), .A1(n35076), .B0(n28326), .C0(n28325), .Y(
        n28359) );
  NAND4XL U32176 ( .A(n28338), .B(n28328), .C(n28327), .D(n28359), .Y(n28361)
         );
  OR2XL U32177 ( .A(n28328), .B(n28327), .Y(n28358) );
  AOI22XL U32178 ( .A0(n34961), .A1(n28330), .B0(n16663), .B1(n28329), .Y(
        n28337) );
  OAI22XL U32179 ( .A0(n28332), .A1(n26621), .B0(n28331), .B1(n16672), .Y(
        n28335) );
  OAI2BB2XL U32180 ( .B0(n35081), .B1(n28333), .A0N(n35079), .A1N(n16670), .Y(
        n28334) );
  AOI211XL U32181 ( .A0(n34827), .A1(n35088), .B0(n28335), .C0(n28334), .Y(
        n28336) );
  OAI211XL U32182 ( .A0(n35085), .A1(n28575), .B0(n28337), .C0(n28336), .Y(
        n28379) );
  INVXL U32183 ( .A(n28338), .Y(n28392) );
  OAI22XL U32184 ( .A0(n35113), .A1(n28575), .B0(n35112), .B1(n18196), .Y(
        n28343) );
  INVXL U32185 ( .A(n28339), .Y(n35117) );
  AOI22XL U32186 ( .A0(n16665), .A1(n35117), .B0(n16663), .B1(n35116), .Y(
        n28341) );
  AOI22XL U32187 ( .A0(n28366), .A1(n35115), .B0(n35114), .B1(n28372), .Y(
        n28340) );
  OAI211XL U32188 ( .A0(n26575), .A1(n35120), .B0(n28341), .C0(n28340), .Y(
        n28342) );
  AOI211XL U32189 ( .A0(n18463), .A1(n35123), .B0(n28343), .C0(n28342), .Y(
        n28380) );
  OAI22XL U32190 ( .A0(n35030), .A1(n28349), .B0(n35033), .B1(n28575), .Y(
        n28348) );
  AOI22XL U32191 ( .A0(n28366), .A1(n35040), .B0(n18463), .B1(n35032), .Y(
        n28346) );
  AOI22XL U32192 ( .A0(n16665), .A1(n28344), .B0(n35034), .B1(n28372), .Y(
        n28345) );
  OAI211XL U32193 ( .A0(n26575), .A1(n35037), .B0(n28346), .C0(n28345), .Y(
        n28347) );
  AOI211XL U32194 ( .A0(n34961), .A1(n35031), .B0(n28348), .C0(n28347), .Y(
        n28381) );
  OAI22XL U32195 ( .A0(n35053), .A1(n28349), .B0(n35055), .B1(n16672), .Y(
        n28356) );
  AOI22XL U32196 ( .A0(n28414), .A1(n28350), .B0(n28366), .B1(n35061), .Y(
        n28354) );
  AOI22XL U32197 ( .A0(n34961), .A1(n28352), .B0(n16670), .B1(n28351), .Y(
        n28353) );
  OAI211XL U32198 ( .A0(n26575), .A1(n35064), .B0(n28354), .C0(n28353), .Y(
        n28355) );
  AOI211XL U32199 ( .A0(n35054), .A1(n28372), .B0(n28356), .C0(n28355), .Y(
        n28385) );
  NAND4XL U32200 ( .A(n28392), .B(n28380), .C(n28381), .D(n28385), .Y(n28357)
         );
  OAI22XL U32201 ( .A0(n28363), .A1(n16672), .B0(n35182), .B1(n18196), .Y(
        n28370) );
  AOI22XL U32202 ( .A0(n28414), .A1(n35185), .B0(n28364), .B1(n28372), .Y(
        n28368) );
  AOI22XL U32203 ( .A0(n28366), .A1(n35179), .B0(n16663), .B1(n28365), .Y(
        n28367) );
  OAI211XL U32204 ( .A0(n26575), .A1(n35192), .B0(n28368), .C0(n28367), .Y(
        n28369) );
  AOI211XL U32205 ( .A0(n16665), .A1(n35189), .B0(n28370), .C0(n28369), .Y(
        n28384) );
  INVXL U32206 ( .A(n28371), .Y(n35203) );
  OAI22XL U32207 ( .A0(n35203), .A1(n16672), .B0(n35201), .B1(n18196), .Y(
        n28378) );
  AOI22XL U32208 ( .A0(n16663), .A1(n28373), .B0(n35206), .B1(n28372), .Y(
        n28376) );
  AOI22XL U32209 ( .A0(n28414), .A1(n28374), .B0(n28366), .B1(n35194), .Y(
        n28375) );
  OAI211XL U32210 ( .A0(n26575), .A1(n35210), .B0(n28376), .C0(n28375), .Y(
        n28377) );
  AOI211XL U32211 ( .A0(n16665), .A1(n35193), .B0(n28378), .C0(n28377), .Y(
        n28383) );
  INVXL U32212 ( .A(pool[109]), .Y(n28393) );
  NAND3XL U32213 ( .A(n28384), .B(n28383), .C(n28393), .Y(n28387) );
  NAND4BBXL U32214 ( .AN(n28381), .BN(n28380), .C(pool[109]), .D(n28379), .Y(
        n28382) );
  AOI22XL U32215 ( .A0(n35010), .A1(n28393), .B0(n28392), .B1(n35006), .Y(
        N29325) );
  OAI2BB1XL U32216 ( .A0N(n28398), .A1N(n28397), .B0(n28396), .Y(n33346) );
  AOI22XL U32217 ( .A0(affine_2[30]), .A1(n33367), .B0(n16674), .B1(n28401), 
        .Y(n28402) );
  NAND2XL U32218 ( .A(n28402), .B(n33350), .Y(n16531) );
  NAND2XL U32219 ( .A(n28404), .B(n28403), .Y(n28409) );
  NAND2XL U32220 ( .A(n28407), .B(n34848), .Y(n28405) );
  OAI211XL U32221 ( .A0(n34851), .A1(n25123), .B0(n28405), .C0(n34831), .Y(
        n34828) );
  AOI22XL U32222 ( .A0(n22362), .A1(n34846), .B0(n28407), .B1(n28406), .Y(
        n28408) );
  NAND2XL U32223 ( .A(n28408), .B(n34831), .Y(n34826) );
  AOI222XL U32224 ( .A0(n28409), .A1(n28467), .B0(n34828), .B1(n28465), .C0(
        n34826), .C1(n26470), .Y(n28598) );
  AOI22XL U32225 ( .A0(n16667), .A1(n28411), .B0(n16660), .B1(n28410), .Y(
        n28424) );
  AOI22XL U32226 ( .A0(n28414), .A1(n28413), .B0(n28559), .B1(n28412), .Y(
        n28423) );
  OAI22XL U32227 ( .A0(n28416), .A1(n28479), .B0(n28415), .B1(n16661), .Y(
        n28420) );
  OAI22XL U32228 ( .A0(n28418), .A1(n28553), .B0(n28417), .B1(n26621), .Y(
        n28419) );
  AOI211XL U32229 ( .A0(n28421), .A1(n28571), .B0(n28420), .C0(n28419), .Y(
        n28422) );
  NAND3XL U32230 ( .A(n28424), .B(n28423), .C(n28422), .Y(n28594) );
  AOI222XL U32231 ( .A0(n28427), .A1(n28467), .B0(n28426), .B1(n28465), .C0(
        n28425), .C1(n35130), .Y(n30644) );
  OAI222XL U32232 ( .A0(n35135), .A1(n28430), .B0(n34989), .B1(n28429), .C0(
        n28428), .C1(N18471), .Y(n34819) );
  AOI222XL U32233 ( .A0(n28433), .A1(n28467), .B0(n28432), .B1(n28465), .C0(
        n28431), .C1(n26470), .Y(n34818) );
  AOI222XL U32234 ( .A0(pool[25]), .A1(pool[26]), .B0(pool[25]), .B1(n34818), 
        .C0(pool[26]), .C1(n34818), .Y(n28434) );
  AOI222XL U32235 ( .A0(n34820), .A1(n34819), .B0(n34820), .B1(n28434), .C0(
        n34819), .C1(n28434), .Y(n28435) );
  AOI222XL U32236 ( .A0(n30644), .A1(pool[28]), .B0(n30644), .B1(n28435), .C0(
        pool[28]), .C1(n28435), .Y(n28548) );
  AOI22XL U32237 ( .A0(n16665), .A1(n28437), .B0(n28571), .B1(n28436), .Y(
        n28448) );
  OAI22XL U32238 ( .A0(n28439), .A1(n28575), .B0(n28438), .B1(n16672), .Y(
        n28446) );
  OAI22XL U32239 ( .A0(n28441), .A1(n16661), .B0(n28440), .B1(n26621), .Y(
        n28445) );
  OAI22XL U32240 ( .A0(n28443), .A1(n28479), .B0(n28442), .B1(n28577), .Y(
        n28444) );
  NOR3XL U32241 ( .A(n28446), .B(n28445), .C(n28444), .Y(n28447) );
  OAI211XL U32242 ( .A0(n28449), .A1(n35198), .B0(n28448), .C0(n28447), .Y(
        n28587) );
  AOI22XL U32243 ( .A0(n28324), .A1(n28451), .B0(n28571), .B1(n28450), .Y(
        n28462) );
  OAI22XL U32244 ( .A0(n28453), .A1(n16661), .B0(n28452), .B1(n28479), .Y(
        n28460) );
  OAI22XL U32245 ( .A0(n28455), .A1(n28575), .B0(n28454), .B1(n28577), .Y(
        n28459) );
  OAI22XL U32246 ( .A0(n28457), .A1(n16672), .B0(n28456), .B1(n28553), .Y(
        n28458) );
  NOR3XL U32247 ( .A(n28460), .B(n28459), .C(n28458), .Y(n28461) );
  OAI211XL U32248 ( .A0(n28463), .A1(n35198), .B0(n28462), .C0(n28461), .Y(
        n28569) );
  AOI222XL U32249 ( .A0(n28468), .A1(n28467), .B0(n28466), .B1(n28465), .C0(
        n28464), .C1(n26470), .Y(n30646) );
  OAI22XL U32250 ( .A0(n28551), .A1(n28470), .B0(n28469), .B1(n16661), .Y(
        n28483) );
  OAI22XL U32251 ( .A0(n28472), .A1(n28553), .B0(n28471), .B1(n28575), .Y(
        n28482) );
  AOI22XL U32252 ( .A0(n16667), .A1(n28474), .B0(n18463), .B1(n28473), .Y(
        n28478) );
  AOI22XL U32253 ( .A0(n18197), .A1(n28476), .B0(n28324), .B1(n28475), .Y(
        n28477) );
  OAI211XL U32254 ( .A0(n28480), .A1(n28479), .B0(n28478), .C0(n28477), .Y(
        n28481) );
  NOR3XL U32255 ( .A(n28483), .B(n28482), .C(n28481), .Y(n28543) );
  AOI22XL U32256 ( .A0(n28528), .A1(n28485), .B0(n28556), .B1(n28484), .Y(
        n28497) );
  AOI22XL U32257 ( .A0(n28366), .A1(n28487), .B0(n28559), .B1(n28486), .Y(
        n28496) );
  OAI22XL U32258 ( .A0(n28489), .A1(n28553), .B0(n28488), .B1(n16661), .Y(
        n28493) );
  OAI22XL U32259 ( .A0(n28491), .A1(n35198), .B0(n28490), .B1(n28575), .Y(
        n28492) );
  AOI211XL U32260 ( .A0(n28571), .A1(n28494), .B0(n28493), .C0(n28492), .Y(
        n28495) );
  NAND3XL U32261 ( .A(n28497), .B(n28496), .C(n28495), .Y(n28545) );
  AOI22XL U32262 ( .A0(n28528), .A1(n28499), .B0(n28324), .B1(n28498), .Y(
        n28510) );
  OAI22XL U32263 ( .A0(n28501), .A1(n16661), .B0(n28500), .B1(n28577), .Y(
        n28508) );
  OAI22XL U32264 ( .A0(n28503), .A1(n35198), .B0(n28502), .B1(n28553), .Y(
        n28507) );
  OAI22XL U32265 ( .A0(n28505), .A1(n16672), .B0(n28504), .B1(n28575), .Y(
        n28506) );
  NOR3XL U32266 ( .A(n28508), .B(n28507), .C(n28506), .Y(n28509) );
  OAI211XL U32267 ( .A0(n28551), .A1(n28511), .B0(n28510), .C0(n28509), .Y(
        n28544) );
  AOI22XL U32268 ( .A0(n16667), .A1(n28513), .B0(n28559), .B1(n28512), .Y(
        n28525) );
  AOI22XL U32269 ( .A0(n16660), .A1(n28515), .B0(n28324), .B1(n28514), .Y(
        n28524) );
  OAI22XL U32270 ( .A0(n28551), .A1(n28517), .B0(n28516), .B1(n16661), .Y(
        n28521) );
  OAI22XL U32271 ( .A0(n28519), .A1(n28553), .B0(n28518), .B1(n28575), .Y(
        n28520) );
  AOI211XL U32272 ( .A0(n34992), .A1(n28522), .B0(n28521), .C0(n28520), .Y(
        n28523) );
  NAND3XL U32273 ( .A(n28525), .B(n28524), .C(n28523), .Y(n28568) );
  AOI22XL U32274 ( .A0(n28528), .A1(n28527), .B0(n16660), .B1(n28526), .Y(
        n28540) );
  AOI22XL U32275 ( .A0(n28366), .A1(n28530), .B0(n28559), .B1(n28529), .Y(
        n28539) );
  OAI22XL U32276 ( .A0(n28532), .A1(n28575), .B0(n28531), .B1(n16661), .Y(
        n28536) );
  OAI22XL U32277 ( .A0(n28551), .A1(n28534), .B0(n28533), .B1(n28553), .Y(
        n28535) );
  AOI211XL U32278 ( .A0(n16667), .A1(n28537), .B0(n28536), .C0(n28535), .Y(
        n28538) );
  NAND3XL U32279 ( .A(n28540), .B(n28539), .C(n28538), .Y(n28567) );
  NOR4XL U32280 ( .A(n28545), .B(n28544), .C(n28568), .D(n28567), .Y(n28541)
         );
  NAND4XL U32281 ( .A(n28542), .B(n30646), .C(n28543), .D(n28541), .Y(n28547)
         );
  OAI22XL U32282 ( .A0(n28551), .A1(n28550), .B0(n28549), .B1(n16661), .Y(
        n28566) );
  OAI22XL U32283 ( .A0(n28554), .A1(n28553), .B0(n28552), .B1(n35198), .Y(
        n28565) );
  AOI22XL U32284 ( .A0(n28528), .A1(n28557), .B0(n28556), .B1(n28555), .Y(
        n28562) );
  AOI22XL U32285 ( .A0(n28324), .A1(n28560), .B0(n28559), .B1(n28558), .Y(
        n28561) );
  OAI211XL U32286 ( .A0(n28563), .A1(n28575), .B0(n28562), .C0(n28561), .Y(
        n28564) );
  OR3XL U32287 ( .A(n28566), .B(n28565), .C(n28564), .Y(n28589) );
  AOI22XL U32288 ( .A0(n16659), .A1(n28572), .B0(n28571), .B1(n28570), .Y(
        n28586) );
  AOI22XL U32289 ( .A0(n18197), .A1(n28574), .B0(n28324), .B1(n28573), .Y(
        n28585) );
  OAI22XL U32290 ( .A0(n28578), .A1(n28577), .B0(n28576), .B1(n28575), .Y(
        n28582) );
  OAI22XL U32291 ( .A0(n28580), .A1(n16661), .B0(n28579), .B1(n16672), .Y(
        n28581) );
  AOI211XL U32292 ( .A0(n16665), .A1(n28583), .B0(n28582), .C0(n28581), .Y(
        n28584) );
  NAND3XL U32293 ( .A(n28586), .B(n28585), .C(n28584), .Y(n28590) );
  NAND4XL U32294 ( .A(pool[29]), .B(n28588), .C(n28590), .D(n28587), .Y(n28592) );
  NOR3XL U32295 ( .A(pool[29]), .B(n28590), .C(n28589), .Y(n28591) );
  NAND2XL U32296 ( .A(n34821), .B(pool[25]), .Y(n28597) );
  OAI21XL U32297 ( .A0(n28598), .A1(n34821), .B0(n28597), .Y(N29241) );
  NAND3XL U32298 ( .A(n34300), .B(conv_1[222]), .C(n28602), .Y(n34678) );
  INVXL U32299 ( .A(conv_1[222]), .Y(n34304) );
  OR2XL U32300 ( .A(n28602), .B(n28601), .Y(n34299) );
  NAND3XL U32301 ( .A(n35392), .B(n34304), .C(n34299), .Y(n34677) );
  AOI22XL U32302 ( .A0(conv_1[223]), .A1(n34678), .B0(n34677), .B1(n34681), 
        .Y(n28604) );
  NAND2XL U32303 ( .A(conv_1[224]), .B(n28604), .Y(n28603) );
  OAI211XL U32304 ( .A0(conv_1[224]), .A1(n28604), .B0(n31735), .C0(n28603), 
        .Y(n28605) );
  OAI211XL U32305 ( .A0(n33853), .A1(n28606), .B0(n16652), .C0(n28605), .Y(
        n16239) );
  OAI2BB1XL U32306 ( .A0N(n28611), .A1N(n28610), .B0(n28609), .Y(n33363) );
  ADDFX1 U32307 ( .A(DP_OP_5171J1_127_4278_n25), .B(n28613), .CI(n28612), .CO(
        n33359), .S(n24575) );
  AOI22XL U32308 ( .A0(affine_2[14]), .A1(n33367), .B0(n16674), .B1(n28614), 
        .Y(n28615) );
  NAND2XL U32309 ( .A(n28615), .B(n33368), .Y(n16565) );
  AOI22XL U32310 ( .A0(n34806), .A1(n28617), .B0(n28616), .B1(n34802), .Y(
        N29230) );
  AOI22XL U32311 ( .A0(n34806), .A1(n28619), .B0(n28618), .B1(n34802), .Y(
        N29229) );
  OAI21XL U32312 ( .A0(n28620), .A1(n16654), .B0(n31191), .Y(n28621) );
  AOI32XL U32313 ( .A0(n34742), .A1(n28621), .A2(n34498), .B0(conv_3[525]), 
        .B1(n28621), .Y(n28622) );
  NAND2XL U32314 ( .A(n34755), .B(n28622), .Y(n15888) );
  INVXL U32315 ( .A(conv_3[148]), .Y(n32169) );
  INVXL U32316 ( .A(conv_3[144]), .Y(n31712) );
  ADDFXL U32317 ( .A(conv_3[142]), .B(n33466), .CI(n28623), .CO(n31720), .S(
        n23779) );
  NAND2XL U32318 ( .A(conv_3[143]), .B(n31720), .Y(n31708) );
  OAI2BB1XL U32319 ( .A0N(conv_3[145]), .A1N(n33465), .B0(n32789), .Y(n33966)
         );
  NAND4XL U32320 ( .A(conv_3[146]), .B(conv_3[147]), .C(n32789), .D(n33966), 
        .Y(n32171) );
  NAND3XL U32321 ( .A(n32788), .B(n33466), .C(n32793), .Y(n32170) );
  NAND2XL U32322 ( .A(n32171), .B(n32170), .Y(n28625) );
  OAI21XL U32323 ( .A0(n16654), .A1(n28625), .B0(n34737), .Y(n28624) );
  AOI32XL U32324 ( .A0(n33778), .A1(n32169), .A2(n28625), .B0(conv_3[148]), 
        .B1(n28624), .Y(n28626) );
  NAND2XL U32325 ( .A(n28626), .B(n35588), .Y(n15645) );
  AOI22XL U32326 ( .A0(n34028), .A1(n28629), .B0(conv_2[312]), .B1(n34026), 
        .Y(n28630) );
  NAND2XL U32327 ( .A(n28630), .B(n35859), .Y(n14996) );
  NAND2XL U32328 ( .A(n34623), .B(n28631), .Y(n28632) );
  INVXL U32329 ( .A(n28632), .Y(n28636) );
  AOI32XL U32330 ( .A0(n34625), .A1(n34631), .A2(n28632), .B0(n36001), .B1(
        n34631), .Y(n28633) );
  AOI21XL U32331 ( .A0(conv_2[159]), .A1(n28633), .B0(n16651), .Y(n28634) );
  OAI31XL U32332 ( .A0(n28636), .A1(n34389), .A2(n28635), .B0(n28634), .Y(
        n15099) );
  ADDFX1 U32333 ( .A(conv_3[10]), .B(n34379), .CI(n28637), .CO(n34378), .S(
        n24374) );
  OAI21XL U32334 ( .A0(conv_3[11]), .A1(n34378), .B0(n34379), .Y(n28639) );
  OAI2BB1XL U32335 ( .A0N(conv_3[11]), .A1N(n34378), .B0(n32996), .Y(n28638)
         );
  AOI31XL U32336 ( .A0(n36020), .A1(n32997), .A2(n28638), .B0(n16653), .Y(
        n28642) );
  OAI2BB1XL U32337 ( .A0N(n28639), .A1N(n28638), .B0(n32656), .Y(n28641) );
  INVXL U32338 ( .A(n28650), .Y(n28645) );
  AOI32XL U32339 ( .A0(n28646), .A1(n33863), .A2(n28645), .B0(n16654), .B1(
        n33863), .Y(n28647) );
  AOI21XL U32340 ( .A0(conv_1[308]), .A1(n28647), .B0(n35549), .Y(n28648) );
  OAI31XL U32341 ( .A0(n28650), .A1(n36042), .A2(n28649), .B0(n28648), .Y(
        n16155) );
  NAND2XL U32342 ( .A(n34706), .B(n29046), .Y(n28654) );
  AOI222XL U32343 ( .A0(n28652), .A1(n28651), .B0(n28652), .B1(conv_2[183]), 
        .C0(n28651), .C1(conv_2[183]), .Y(n28653) );
  NOR2X1 U32344 ( .A(conv_2[189]), .B(n28657), .Y(n29891) );
  NAND2XL U32345 ( .A(conv_2[186]), .B(n29910), .Y(n29886) );
  NAND2XL U32346 ( .A(conv_2[188]), .B(n35913), .Y(n29892) );
  NAND2XL U32347 ( .A(n30946), .B(n29892), .Y(n28656) );
  AOI32XL U32348 ( .A0(n29892), .A1(n36020), .A2(n30946), .B0(n28657), .B1(
        n36020), .Y(n28658) );
  AOI32XL U32349 ( .A0(n35917), .A1(n28659), .A2(n28658), .B0(n29893), .B1(
        n28659), .Y(n15079) );
  INVXL U32350 ( .A(n33770), .Y(n31121) );
  NAND2XL U32351 ( .A(n31121), .B(n30428), .Y(n28666) );
  AOI32XL U32352 ( .A0(n30428), .A1(n36020), .A2(n31121), .B0(n28667), .B1(
        n36020), .Y(n28668) );
  AOI32XL U32353 ( .A0(n35934), .A1(n28669), .A2(n28668), .B0(n30429), .B1(
        n28669), .Y(n15059) );
  NAND2XL U32354 ( .A(n28673), .B(n28674), .Y(n28670) );
  AOI32XL U32355 ( .A0(n28674), .A1(n36020), .A2(n28673), .B0(n28672), .B1(
        n33157), .Y(n28676) );
  AOI32XL U32356 ( .A0(n30412), .A1(n28677), .A2(n28676), .B0(n28675), .B1(
        n28677), .Y(n15189) );
  NAND2XL U32357 ( .A(n28679), .B(n28678), .Y(n30143) );
  INVXL U32358 ( .A(conv_2[112]), .Y(n35886) );
  OAI2BB1XL U32359 ( .A0N(conv_2[110]), .A1N(n28680), .B0(n35884), .Y(n30142)
         );
  NAND2XL U32360 ( .A(conv_2[111]), .B(n30142), .Y(n35883) );
  NAND2XL U32361 ( .A(conv_2[113]), .B(n35890), .Y(n30135) );
  NAND2XL U32362 ( .A(n35884), .B(n30135), .Y(n28681) );
  AOI32XL U32363 ( .A0(n30135), .A1(n36020), .A2(n35884), .B0(n28682), .B1(
        n33778), .Y(n28683) );
  AOI32XL U32364 ( .A0(n35894), .A1(n28684), .A2(n28683), .B0(n30136), .B1(
        n28684), .Y(n15129) );
  AOI22XL U32365 ( .A0(conv_3[5]), .A1(n34379), .B0(n32996), .B1(n28689), .Y(
        n28686) );
  NAND2XL U32366 ( .A(n28687), .B(n28686), .Y(n28685) );
  OAI211XL U32367 ( .A0(n28687), .A1(n28686), .B0(n33157), .C0(n28685), .Y(
        n28688) );
  OAI211XL U32368 ( .A0(n34383), .A1(n28689), .B0(n16649), .C0(n28688), .Y(
        n15743) );
  INVXL U32369 ( .A(n28691), .Y(n28695) );
  AOI32XL U32370 ( .A0(n28691), .A1(n34447), .A2(n28690), .B0(n16655), .B1(
        n34447), .Y(n28692) );
  AOI21XL U32371 ( .A0(conv_2[95]), .A1(n28692), .B0(n16651), .Y(n28693) );
  OAI31XL U32372 ( .A0(n28695), .A1(n36042), .A2(n28694), .B0(n28693), .Y(
        n15143) );
  NAND2XL U32373 ( .A(n30225), .B(n28696), .Y(n28697) );
  INVXL U32374 ( .A(n28697), .Y(n28702) );
  AOI32XL U32375 ( .A0(n28698), .A1(n34447), .A2(n28697), .B0(n16654), .B1(
        n34447), .Y(n28699) );
  AOI21XL U32376 ( .A0(conv_2[96]), .A1(n28699), .B0(n16651), .Y(n28700) );
  OAI31XL U32377 ( .A0(n28702), .A1(n36042), .A2(n28701), .B0(n28700), .Y(
        n15142) );
  NAND2XL U32378 ( .A(n28706), .B(n28707), .Y(n28703) );
  AOI31XL U32379 ( .A0(n16657), .A1(n28704), .A2(n28703), .B0(n16651), .Y(
        n28710) );
  AOI32XL U32380 ( .A0(n28707), .A1(n36020), .A2(n28706), .B0(n28705), .B1(
        n33157), .Y(n28709) );
  NAND2XL U32381 ( .A(n31134), .B(n28714), .Y(n28711) );
  AOI31XL U32382 ( .A0(n16656), .A1(n28712), .A2(n28711), .B0(n16651), .Y(
        n28717) );
  AOI32XL U32383 ( .A0(n28714), .A1(n36020), .A2(n31134), .B0(n28713), .B1(
        n16657), .Y(n28716) );
  AOI32XL U32384 ( .A0(n34505), .A1(n28717), .A2(n28716), .B0(n28715), .B1(
        n28717), .Y(n15169) );
  OAI21XL U32385 ( .A0(n28718), .A1(n16654), .B0(n35805), .Y(n28719) );
  AOI32XL U32386 ( .A0(n34742), .A1(n28719), .A2(n34444), .B0(conv_3[450]), 
        .B1(n28719), .Y(n28720) );
  NAND2XL U32387 ( .A(n34755), .B(n28720), .Y(n15893) );
  NAND2XL U32388 ( .A(n33478), .B(n28724), .Y(n29113) );
  NAND2XL U32389 ( .A(conv_3[260]), .B(n29113), .Y(n29131) );
  NAND2XL U32390 ( .A(n29107), .B(conv_3[262]), .Y(n32101) );
  NAND2XL U32391 ( .A(n33478), .B(n32101), .Y(n28725) );
  AOI31XL U32392 ( .A0(n16657), .A1(n32102), .A2(n28725), .B0(n16653), .Y(
        n28728) );
  AOI32XL U32393 ( .A0(n32101), .A1(n36020), .A2(n33478), .B0(n28726), .B1(
        n36020), .Y(n28727) );
  AOI32XL U32394 ( .A0(n35713), .A1(n28728), .A2(n28727), .B0(n32100), .B1(
        n28728), .Y(n15570) );
  NAND3XL U32395 ( .A(conv_1[462]), .B(n30051), .C(n28729), .Y(n28749) );
  NAND3XL U32396 ( .A(n30044), .B(n28731), .C(n28730), .Y(n28748) );
  NAND2XL U32397 ( .A(n28749), .B(n28748), .Y(n28733) );
  NAND2XL U32398 ( .A(conv_1[463]), .B(n28733), .Y(n28732) );
  OAI211XL U32399 ( .A0(conv_1[463]), .A1(n28733), .B0(n28751), .C0(n28732), 
        .Y(n28734) );
  OAI211XL U32400 ( .A0(n30056), .A1(n28747), .B0(n34689), .C0(n28734), .Y(
        n16000) );
  INVXL U32401 ( .A(weight_1[215]), .Y(n32912) );
  INVXL U32402 ( .A(weight_1[221]), .Y(n32816) );
  OAI22XL U32403 ( .A0(n16645), .A1(n32912), .B0(n32816), .B1(n16647), .Y(
        n14141) );
  INVXL U32404 ( .A(weight_1[287]), .Y(n32802) );
  INVXL U32405 ( .A(weight_1[293]), .Y(n32800) );
  OAI22XL U32406 ( .A0(n32491), .A1(n32802), .B0(n32800), .B1(n26910), .Y(
        n14153) );
  INVXL U32407 ( .A(weight_1[251]), .Y(n32807) );
  INVXL U32408 ( .A(weight_1[257]), .Y(n32801) );
  OAI22XL U32409 ( .A0(n31084), .A1(n32807), .B0(n32801), .B1(n16647), .Y(
        n14147) );
  NAND4XL U32410 ( .A(conv_1[476]), .B(conv_1[477]), .C(n29824), .D(n29823), 
        .Y(n33245) );
  NAND3XL U32411 ( .A(n32887), .B(n29821), .C(n29828), .Y(n33244) );
  AOI22XL U32412 ( .A0(conv_1[478]), .A1(n33245), .B0(n33244), .B1(n33248), 
        .Y(n28736) );
  NAND2XL U32413 ( .A(conv_1[479]), .B(n28736), .Y(n28735) );
  OAI211XL U32414 ( .A0(conv_1[479]), .A1(n28736), .B0(n32181), .C0(n28735), 
        .Y(n28737) );
  OAI211XL U32415 ( .A0(n33853), .A1(n28738), .B0(n16652), .C0(n28737), .Y(
        n15984) );
  INVXL U32416 ( .A(conv_2[82]), .Y(n30171) );
  NAND2XL U32417 ( .A(conv_2[81]), .B(n35869), .Y(n30167) );
  NAND2XL U32418 ( .A(conv_2[83]), .B(n35875), .Y(n30173) );
  NAND2XL U32419 ( .A(n30924), .B(n30173), .Y(n28743) );
  AOI31XL U32420 ( .A0(n36020), .A1(n30172), .A2(n28743), .B0(n16651), .Y(
        n28746) );
  AOI32XL U32421 ( .A0(n30173), .A1(n36020), .A2(n30924), .B0(n28744), .B1(
        n16657), .Y(n28745) );
  AOI22XL U32422 ( .A0(conv_1[463]), .A1(n28749), .B0(n28748), .B1(n28747), 
        .Y(n28752) );
  NAND2XL U32423 ( .A(conv_1[464]), .B(n28752), .Y(n28750) );
  OAI211XL U32424 ( .A0(conv_1[464]), .A1(n28752), .B0(n28751), .C0(n28750), 
        .Y(n28753) );
  OAI211XL U32425 ( .A0(n33442), .A1(n28754), .B0(n34689), .C0(n28753), .Y(
        n15999) );
  NOR2X1 U32426 ( .A(n33281), .B(n28757), .Y(n31901) );
  NAND2XL U32427 ( .A(n33281), .B(n28757), .Y(n31902) );
  NAND2XL U32428 ( .A(n33281), .B(n31909), .Y(n28758) );
  AOI31XL U32429 ( .A0(n36020), .A1(n31907), .A2(n28758), .B0(n16653), .Y(
        n28761) );
  AOI32XL U32430 ( .A0(n31909), .A1(n36020), .A2(n33281), .B0(n28759), .B1(
        n36020), .Y(n28760) );
  INVXL U32431 ( .A(conv_3[321]), .Y(n31908) );
  INVXL U32432 ( .A(conv_3[165]), .Y(n28764) );
  OAI2BB1XL U32433 ( .A0N(n36020), .A1N(n28762), .B0(n35630), .Y(n28763) );
  AOI32XL U32434 ( .A0(n34742), .A1(n28764), .A2(n34433), .B0(conv_3[165]), 
        .B1(n28763), .Y(n28765) );
  NAND2XL U32435 ( .A(n28765), .B(n34755), .Y(n15912) );
  OAI21XL U32436 ( .A0(n35950), .A1(n28767), .B0(n28766), .Y(n28769) );
  AOI211XL U32437 ( .A0(n28771), .A1(n28769), .B0(n36042), .C0(n28768), .Y(
        n28770) );
  AOI2BB1XL U32438 ( .A0N(n28771), .A1N(n30994), .B0(n28770), .Y(n28772) );
  NAND2XL U32439 ( .A(n35859), .B(n28772), .Y(n15021) );
  INVXL U32440 ( .A(conv_2[5]), .Y(n30959) );
  NAND2XL U32441 ( .A(n33571), .B(intadd_0_n1), .Y(n30954) );
  AOI32XL U32442 ( .A0(n30959), .A1(n28773), .A2(n30954), .B0(n29583), .B1(
        n28773), .Y(n28775) );
  NAND2XL U32443 ( .A(n28777), .B(n28775), .Y(n28774) );
  OAI211XL U32444 ( .A0(n28777), .A1(n28775), .B0(n33788), .C0(n28774), .Y(
        n28776) );
  OAI211XL U32445 ( .A0(n30958), .A1(n28777), .B0(n34669), .C0(n28776), .Y(
        n15202) );
  AOI21XL U32446 ( .A0(n29583), .A1(n28779), .B0(n28778), .Y(n28781) );
  NAND2XL U32447 ( .A(conv_2[9]), .B(n28781), .Y(n28780) );
  OAI211XL U32448 ( .A0(conv_2[9]), .A1(n28781), .B0(n36020), .C0(n28780), .Y(
        n28782) );
  OAI211XL U32449 ( .A0(n30958), .A1(n28783), .B0(n33815), .C0(n28782), .Y(
        n15199) );
  AOI2BB1XL U32450 ( .A0N(n33571), .A1N(n28785), .B0(n28784), .Y(n28787) );
  NAND2XL U32451 ( .A(conv_2[10]), .B(n28787), .Y(n28786) );
  OAI211XL U32452 ( .A0(conv_2[10]), .A1(n28787), .B0(n36020), .C0(n28786), 
        .Y(n28788) );
  OAI211XL U32453 ( .A0(n30958), .A1(n28789), .B0(n35859), .C0(n28788), .Y(
        n15198) );
  AOI21XL U32454 ( .A0(n28937), .A1(n28791), .B0(n28790), .Y(n28793) );
  NAND2XL U32455 ( .A(conv_2[444]), .B(n28793), .Y(n28792) );
  OAI211XL U32456 ( .A0(conv_2[444]), .A1(n28793), .B0(n32656), .C0(n28792), 
        .Y(n28794) );
  OAI211XL U32457 ( .A0(n36070), .A1(n28795), .B0(n34669), .C0(n28794), .Y(
        n14909) );
  NAND2XL U32458 ( .A(conv_3[246]), .B(n35680), .Y(n35686) );
  NAND2XL U32459 ( .A(conv_3[248]), .B(n35692), .Y(n35699) );
  AOI221XL U32460 ( .A0(n28800), .A1(n16656), .B0(n28799), .B1(n33788), .C0(
        n33545), .Y(n28803) );
  INVXL U32461 ( .A(conv_3[250]), .Y(n28802) );
  OAI211XL U32462 ( .A0(n35693), .A1(n29118), .B0(n33822), .C0(n29119), .Y(
        n28801) );
  OAI211XL U32463 ( .A0(n28803), .A1(n28802), .B0(n33468), .C0(n28801), .Y(
        n15578) );
  AOI2BB1XL U32464 ( .A0N(n35441), .A1N(n28815), .B0(n28816), .Y(n28806) );
  NAND2XL U32465 ( .A(conv_1[355]), .B(n28806), .Y(n28805) );
  OAI211XL U32466 ( .A0(conv_1[355]), .A1(n28806), .B0(n32611), .C0(n28805), 
        .Y(n28807) );
  OAI211XL U32467 ( .A0(n35447), .A1(n28808), .B0(n16652), .C0(n28807), .Y(
        n16108) );
  NAND2XL U32468 ( .A(conv_1[352]), .B(n28812), .Y(n28811) );
  OAI211XL U32469 ( .A0(conv_1[352]), .A1(n28812), .B0(n32660), .C0(n28811), 
        .Y(n28813) );
  OAI211XL U32470 ( .A0(n35447), .A1(n28814), .B0(n34281), .C0(n28813), .Y(
        n16111) );
  NAND4XL U32471 ( .A(conv_1[356]), .B(conv_1[357]), .C(n28847), .D(n35449), 
        .Y(n33998) );
  OAI21XL U32472 ( .A0(conv_1[355]), .A1(n28816), .B0(n35441), .Y(n35448) );
  INVXL U32473 ( .A(conv_1[357]), .Y(n28851) );
  NAND3XL U32474 ( .A(n35450), .B(n35441), .C(n28851), .Y(n33997) );
  INVXL U32475 ( .A(conv_1[358]), .Y(n34001) );
  AOI22XL U32476 ( .A0(conv_1[358]), .A1(n33998), .B0(n33997), .B1(n34001), 
        .Y(n28818) );
  NAND2XL U32477 ( .A(conv_1[359]), .B(n28818), .Y(n28817) );
  OAI211XL U32478 ( .A0(conv_1[359]), .A1(n28818), .B0(n33157), .C0(n28817), 
        .Y(n28819) );
  OAI211XL U32479 ( .A0(n33442), .A1(n28820), .B0(n16652), .C0(n28819), .Y(
        n16104) );
  NAND4XL U32480 ( .A(conv_1[341]), .B(conv_1[342]), .C(n28821), .D(n33884), 
        .Y(n28842) );
  INVXL U32481 ( .A(conv_1[342]), .Y(n33889) );
  NAND2XL U32482 ( .A(n28823), .B(n28822), .Y(n28824) );
  NAND2XL U32483 ( .A(n35434), .B(n28824), .Y(n33885) );
  NAND3XL U32484 ( .A(n35434), .B(n33889), .C(n33885), .Y(n28841) );
  INVXL U32485 ( .A(conv_1[343]), .Y(n28846) );
  AOI22XL U32486 ( .A0(conv_1[343]), .A1(n28842), .B0(n28841), .B1(n28846), 
        .Y(n28826) );
  NAND2XL U32487 ( .A(conv_1[344]), .B(n28826), .Y(n28825) );
  OAI211XL U32488 ( .A0(conv_1[344]), .A1(n28826), .B0(n33778), .C0(n28825), 
        .Y(n28827) );
  OAI211XL U32489 ( .A0(n33442), .A1(n28828), .B0(n34696), .C0(n28827), .Y(
        n16119) );
  NAND2XL U32490 ( .A(conv_3[216]), .B(n35659), .Y(n31529) );
  NAND2XL U32491 ( .A(n34649), .B(n31529), .Y(n28832) );
  INVXL U32492 ( .A(conv_3[217]), .Y(n31530) );
  NAND2XL U32493 ( .A(conv_3[203]), .B(n34656), .Y(n31846) );
  NAND2XL U32494 ( .A(n31848), .B(n31846), .Y(n28837) );
  AOI32XL U32495 ( .A0(n31846), .A1(n36020), .A2(n31848), .B0(n28838), .B1(
        n36020), .Y(n28839) );
  NAND2XL U32496 ( .A(n28842), .B(n28841), .Y(n28844) );
  NAND2XL U32497 ( .A(conv_1[343]), .B(n28844), .Y(n28843) );
  OAI211XL U32498 ( .A0(conv_1[343]), .A1(n28844), .B0(n16657), .C0(n28843), 
        .Y(n28845) );
  OAI211XL U32499 ( .A0(n35437), .A1(n28846), .B0(n34682), .C0(n28845), .Y(
        n16120) );
  AOI32XL U32500 ( .A0(conv_1[356]), .A1(n28847), .A2(n35449), .B0(n35441), 
        .B1(n35450), .Y(n28849) );
  NAND2XL U32501 ( .A(n28851), .B(n28849), .Y(n28848) );
  OAI211XL U32502 ( .A0(n28851), .A1(n28849), .B0(n34028), .C0(n28848), .Y(
        n28850) );
  OAI211XL U32503 ( .A0(n35447), .A1(n28851), .B0(n34689), .C0(n28850), .Y(
        n16106) );
  INVXL U32504 ( .A(conv_2[529]), .Y(n28857) );
  NAND2XL U32505 ( .A(conv_2[529]), .B(n28855), .Y(n28854) );
  OAI211XL U32506 ( .A0(conv_2[529]), .A1(n28855), .B0(n33778), .C0(n28854), 
        .Y(n28856) );
  OAI211XL U32507 ( .A0(n34496), .A1(n28857), .B0(n28856), .C0(n34408), .Y(
        n15204) );
  NOR2BXL U32508 ( .AN(n28859), .B(n28858), .Y(n28861) );
  NAND2XL U32509 ( .A(conv_2[409]), .B(n28861), .Y(n28860) );
  OAI211XL U32510 ( .A0(conv_2[409]), .A1(n28861), .B0(n16657), .C0(n28860), 
        .Y(n28862) );
  OAI211XL U32511 ( .A0(n36047), .A1(n28863), .B0(n28862), .C0(n34408), .Y(
        n15212) );
  INVXL U32512 ( .A(conv_2[319]), .Y(n28869) );
  NAND2XL U32513 ( .A(conv_2[319]), .B(n28867), .Y(n28866) );
  OAI211XL U32514 ( .A0(conv_2[319]), .A1(n28867), .B0(n36020), .C0(n28866), 
        .Y(n28868) );
  OAI211XL U32515 ( .A0(n35986), .A1(n28869), .B0(n28868), .C0(n34408), .Y(
        n15218) );
  INVXL U32516 ( .A(conv_2[304]), .Y(n28875) );
  NAND2XL U32517 ( .A(conv_2[304]), .B(n28873), .Y(n28872) );
  OAI211XL U32518 ( .A0(conv_2[304]), .A1(n28873), .B0(n33822), .C0(n28872), 
        .Y(n28874) );
  OAI211XL U32519 ( .A0(n35976), .A1(n28875), .B0(n28874), .C0(n34408), .Y(
        n15219) );
  NAND2XL U32520 ( .A(conv_2[214]), .B(n28879), .Y(n28878) );
  OAI211XL U32521 ( .A0(conv_2[214]), .A1(n28879), .B0(n36020), .C0(n28878), 
        .Y(n28880) );
  OAI211XL U32522 ( .A0(n35934), .A1(n28881), .B0(n28880), .C0(n34408), .Y(
        n15225) );
  AOI22XL U32523 ( .A0(n33788), .A1(intadd_1_SUM_2_), .B0(conv_1[425]), .B1(
        n35510), .Y(n28882) );
  NAND2XL U32524 ( .A(n28882), .B(n34689), .Y(n16038) );
  NAND4XL U32525 ( .A(conv_2[281]), .B(conv_2[282]), .C(n28883), .D(n30985), 
        .Y(n30993) );
  INVXL U32526 ( .A(conv_2[282]), .Y(n30990) );
  NAND2XL U32527 ( .A(n28885), .B(n28884), .Y(n28886) );
  NAND2XL U32528 ( .A(n35950), .B(n28886), .Y(n30986) );
  NAND3XL U32529 ( .A(n35950), .B(n30990), .C(n30986), .Y(n30992) );
  INVXL U32530 ( .A(conv_2[283]), .Y(n30997) );
  AOI22XL U32531 ( .A0(conv_2[283]), .A1(n30993), .B0(n30992), .B1(n30997), 
        .Y(n28888) );
  NAND2XL U32532 ( .A(conv_2[284]), .B(n28888), .Y(n28887) );
  OAI211XL U32533 ( .A0(conv_2[284]), .A1(n28888), .B0(n33778), .C0(n28887), 
        .Y(n28889) );
  OAI211XL U32534 ( .A0(n33442), .A1(n28890), .B0(n34735), .C0(n28889), .Y(
        n15014) );
  NAND2XL U32535 ( .A(n28930), .B(conv_2[426]), .Y(n28905) );
  INVXL U32536 ( .A(n34211), .Y(n28906) );
  OAI2BB1XL U32537 ( .A0N(n28924), .A1N(conv_2[428]), .B0(n28906), .Y(n36054)
         );
  OAI21XL U32538 ( .A0(conv_2[428]), .A1(n28923), .B0(n34211), .Y(n36052) );
  NAND4XL U32539 ( .A(conv_2[431]), .B(conv_2[432]), .C(n34210), .D(n28906), 
        .Y(n28912) );
  AOI22XL U32540 ( .A0(conv_2[433]), .A1(n28912), .B0(n28911), .B1(n28916), 
        .Y(n28895) );
  NAND2XL U32541 ( .A(conv_2[434]), .B(n28895), .Y(n28894) );
  OAI211XL U32542 ( .A0(conv_2[434]), .A1(n28895), .B0(n33982), .C0(n28894), 
        .Y(n28896) );
  OAI211XL U32543 ( .A0(n33853), .A1(n28897), .B0(n34669), .C0(n28896), .Y(
        n14914) );
  AOI21XL U32544 ( .A0(n35970), .A1(n28899), .B0(n28898), .Y(n28901) );
  NAND2XL U32545 ( .A(conv_2[307]), .B(n28901), .Y(n28900) );
  OAI211XL U32546 ( .A0(conv_2[307]), .A1(n28901), .B0(n36020), .C0(n28900), 
        .Y(n28902) );
  OAI211XL U32547 ( .A0(n35976), .A1(n28903), .B0(n35859), .C0(n28902), .Y(
        n15001) );
  AOI21XL U32548 ( .A0(n28906), .A1(n28905), .B0(n28904), .Y(n28908) );
  NAND2XL U32549 ( .A(conv_2[427]), .B(n28908), .Y(n28907) );
  OAI211XL U32550 ( .A0(conv_2[427]), .A1(n28908), .B0(n33788), .C0(n28907), 
        .Y(n28909) );
  OAI211XL U32551 ( .A0(n36053), .A1(n28910), .B0(n34735), .C0(n28909), .Y(
        n14921) );
  NAND2XL U32552 ( .A(n28912), .B(n28911), .Y(n28914) );
  NAND2XL U32553 ( .A(conv_2[433]), .B(n28914), .Y(n28913) );
  OAI211XL U32554 ( .A0(conv_2[433]), .A1(n28914), .B0(n16657), .C0(n28913), 
        .Y(n28915) );
  OAI211XL U32555 ( .A0(n36053), .A1(n28916), .B0(n34669), .C0(n28915), .Y(
        n14915) );
  INVXL U32556 ( .A(conv_2[306]), .Y(n28922) );
  AOI2BB1XL U32557 ( .A0N(n33979), .A1N(n28918), .B0(n28917), .Y(n28920) );
  NAND2XL U32558 ( .A(conv_2[306]), .B(n28920), .Y(n28919) );
  OAI211XL U32559 ( .A0(conv_2[306]), .A1(n28920), .B0(n33982), .C0(n28919), 
        .Y(n28921) );
  OAI211XL U32560 ( .A0(n35976), .A1(n28922), .B0(n35859), .C0(n28921), .Y(
        n15002) );
  AOI2BB1XL U32561 ( .A0N(n34211), .A1N(n28924), .B0(n28923), .Y(n28926) );
  NAND2XL U32562 ( .A(conv_2[428]), .B(n28926), .Y(n28925) );
  OAI211XL U32563 ( .A0(conv_2[428]), .A1(n28926), .B0(n16656), .C0(n28925), 
        .Y(n28927) );
  OAI211XL U32564 ( .A0(n36053), .A1(n28928), .B0(n34735), .C0(n28927), .Y(
        n14920) );
  AOI2BB1XL U32565 ( .A0N(n34211), .A1N(n28930), .B0(n28929), .Y(n28932) );
  NAND2XL U32566 ( .A(conv_2[426]), .B(n28932), .Y(n28931) );
  OAI211XL U32567 ( .A0(conv_2[426]), .A1(n28932), .B0(n16657), .C0(n28931), 
        .Y(n28933) );
  OAI211XL U32568 ( .A0(n36053), .A1(n28934), .B0(n34669), .C0(n28933), .Y(
        n14922) );
  AOI21XL U32569 ( .A0(n28937), .A1(n28936), .B0(n28935), .Y(n28939) );
  NAND2XL U32570 ( .A(conv_2[442]), .B(n28939), .Y(n28938) );
  OAI211XL U32571 ( .A0(conv_2[442]), .A1(n28939), .B0(n33788), .C0(n28938), 
        .Y(n28940) );
  OAI211XL U32572 ( .A0(n36070), .A1(n28941), .B0(n34735), .C0(n28940), .Y(
        n14911) );
  NAND2XL U32573 ( .A(conv_2[440]), .B(n28945), .Y(n28944) );
  OAI211XL U32574 ( .A0(conv_2[440]), .A1(n28945), .B0(n30090), .C0(n28944), 
        .Y(n28946) );
  OAI211XL U32575 ( .A0(n36070), .A1(n28947), .B0(n34669), .C0(n28946), .Y(
        n14913) );
  NOR2X1 U32576 ( .A(n35622), .B(n28951), .Y(n31399) );
  AOI2BB1XL U32577 ( .A0N(n35623), .A1N(conv_3[127]), .B0(n34783), .Y(n31412)
         );
  INVXL U32578 ( .A(conv_3[127]), .Y(n35625) );
  NAND2XL U32579 ( .A(n31413), .B(conv_3[128]), .Y(n31437) );
  NAND2XL U32580 ( .A(n34783), .B(n31437), .Y(n28952) );
  AOI31XL U32581 ( .A0(n33712), .A1(n31438), .A2(n28952), .B0(n16653), .Y(
        n28955) );
  AOI32XL U32582 ( .A0(n31437), .A1(n36020), .A2(n34783), .B0(n28953), .B1(
        n16657), .Y(n28954) );
  INVXL U32583 ( .A(conv_3[129]), .Y(n31436) );
  NAND2XL U32584 ( .A(n28959), .B(n28960), .Y(n28956) );
  AOI31XL U32585 ( .A0(n36020), .A1(n28957), .A2(n28956), .B0(n16653), .Y(
        n28963) );
  AOI32XL U32586 ( .A0(n28960), .A1(n36020), .A2(n28959), .B0(n28958), .B1(
        n33778), .Y(n28962) );
  INVXL U32587 ( .A(conv_1[363]), .Y(n28970) );
  AOI21XL U32588 ( .A0(n28966), .A1(n28965), .B0(n28964), .Y(n28968) );
  NAND2XL U32589 ( .A(conv_1[363]), .B(n28968), .Y(n28967) );
  OAI211XL U32590 ( .A0(conv_1[363]), .A1(n28968), .B0(n33788), .C0(n28967), 
        .Y(n28969) );
  OAI211XL U32591 ( .A0(n35458), .A1(n28970), .B0(n32867), .C0(n28969), .Y(
        n16100) );
  INVXL U32592 ( .A(conv_2[514]), .Y(n28976) );
  NAND2XL U32593 ( .A(conv_2[514]), .B(n28974), .Y(n28973) );
  OAI211XL U32594 ( .A0(conv_2[514]), .A1(n28974), .B0(n32611), .C0(n28973), 
        .Y(n28975) );
  OAI211XL U32595 ( .A0(n31013), .A1(n28976), .B0(n34408), .C0(n28975), .Y(
        n15205) );
  NOR2BXL U32596 ( .AN(n28978), .B(n28977), .Y(n28980) );
  NAND2XL U32597 ( .A(conv_2[244]), .B(n28980), .Y(n28979) );
  OAI211XL U32598 ( .A0(conv_2[244]), .A1(n28980), .B0(n36020), .C0(n28979), 
        .Y(n28981) );
  OAI211XL U32599 ( .A0(n35945), .A1(n28982), .B0(n34408), .C0(n28981), .Y(
        n15223) );
  INVXL U32600 ( .A(conv_2[484]), .Y(n28988) );
  NAND2XL U32601 ( .A(conv_2[484]), .B(n28986), .Y(n28985) );
  OAI211XL U32602 ( .A0(conv_2[484]), .A1(n28986), .B0(n32656), .C0(n28985), 
        .Y(n28987) );
  OAI211XL U32603 ( .A0(n34137), .A1(n28988), .B0(n34408), .C0(n28987), .Y(
        n15207) );
  INVXL U32604 ( .A(conv_2[499]), .Y(n28994) );
  NAND2XL U32605 ( .A(conv_2[499]), .B(n28992), .Y(n28991) );
  OAI211XL U32606 ( .A0(conv_2[499]), .A1(n28992), .B0(n33157), .C0(n28991), 
        .Y(n28993) );
  OAI211XL U32607 ( .A0(n36091), .A1(n28994), .B0(n34408), .C0(n28993), .Y(
        n15206) );
  INVXL U32608 ( .A(conv_2[469]), .Y(n29000) );
  NOR2BXL U32609 ( .AN(n28996), .B(n28995), .Y(n28998) );
  NAND2XL U32610 ( .A(conv_2[469]), .B(n28998), .Y(n28997) );
  OAI211XL U32611 ( .A0(conv_2[469]), .A1(n28998), .B0(n33778), .C0(n28997), 
        .Y(n28999) );
  OAI211XL U32612 ( .A0(n34177), .A1(n29000), .B0(n34408), .C0(n28999), .Y(
        n15208) );
  INVXL U32613 ( .A(conv_2[169]), .Y(n29009) );
  INVXL U32614 ( .A(n29003), .Y(n29005) );
  NAND2XL U32615 ( .A(conv_2[169]), .B(n29007), .Y(n29006) );
  OAI211XL U32616 ( .A0(conv_2[169]), .A1(n29007), .B0(n33788), .C0(n29006), 
        .Y(n29008) );
  OAI211XL U32617 ( .A0(n34589), .A1(n29009), .B0(n34408), .C0(n29008), .Y(
        n15228) );
  INVXL U32618 ( .A(conv_2[379]), .Y(n29015) );
  NAND2XL U32619 ( .A(conv_2[379]), .B(n29013), .Y(n29012) );
  OAI211XL U32620 ( .A0(conv_2[379]), .A1(n29013), .B0(n33982), .C0(n29012), 
        .Y(n29014) );
  OAI211XL U32621 ( .A0(n36028), .A1(n29015), .B0(n34408), .C0(n29014), .Y(
        n15214) );
  NAND2XL U32622 ( .A(conv_2[424]), .B(n29019), .Y(n29018) );
  OAI211XL U32623 ( .A0(conv_2[424]), .A1(n29019), .B0(n33778), .C0(n29018), 
        .Y(n29020) );
  OAI211XL U32624 ( .A0(n36053), .A1(n29021), .B0(n34408), .C0(n29020), .Y(
        n15211) );
  INVXL U32625 ( .A(conv_2[184]), .Y(n29027) );
  NAND2XL U32626 ( .A(conv_2[184]), .B(n29025), .Y(n29024) );
  OAI211XL U32627 ( .A0(conv_2[184]), .A1(n29025), .B0(n33982), .C0(n29024), 
        .Y(n29026) );
  OAI211XL U32628 ( .A0(n35917), .A1(n29027), .B0(n34408), .C0(n29026), .Y(
        n15227) );
  NAND2XL U32629 ( .A(conv_2[439]), .B(n29031), .Y(n29030) );
  OAI211XL U32630 ( .A0(conv_2[439]), .A1(n29031), .B0(n16657), .C0(n29030), 
        .Y(n29032) );
  OAI211XL U32631 ( .A0(n36070), .A1(n29033), .B0(n34408), .C0(n29032), .Y(
        n15210) );
  INVXL U32632 ( .A(conv_2[289]), .Y(n29039) );
  NAND2XL U32633 ( .A(conv_2[289]), .B(n29037), .Y(n29036) );
  OAI211XL U32634 ( .A0(conv_2[289]), .A1(n29037), .B0(n36020), .C0(n29036), 
        .Y(n29038) );
  OAI211XL U32635 ( .A0(n35963), .A1(n29039), .B0(n34408), .C0(n29038), .Y(
        n15220) );
  INVXL U32636 ( .A(conv_2[199]), .Y(n29045) );
  NOR2BXL U32637 ( .AN(n29041), .B(n29040), .Y(n29043) );
  NAND2XL U32638 ( .A(conv_2[199]), .B(n29043), .Y(n29042) );
  OAI211XL U32639 ( .A0(conv_2[199]), .A1(n29043), .B0(n36020), .C0(n29042), 
        .Y(n29044) );
  OAI211XL U32640 ( .A0(n35931), .A1(n29045), .B0(n34408), .C0(n29044), .Y(
        n15226) );
  NAND2XL U32641 ( .A(n34461), .B(n29046), .Y(n29050) );
  AOI222XL U32642 ( .A0(n29048), .A1(conv_2[228]), .B0(n29048), .B1(n29047), 
        .C0(conv_2[228]), .C1(n29047), .Y(n29049) );
  NAND2XL U32643 ( .A(n29050), .B(n29049), .Y(n29137) );
  NOR2BXL U32644 ( .AN(n29137), .B(n29138), .Y(n29052) );
  NAND2XL U32645 ( .A(conv_2[229]), .B(n29052), .Y(n29051) );
  OAI211XL U32646 ( .A0(conv_2[229]), .A1(n29052), .B0(n36020), .C0(n29051), 
        .Y(n29053) );
  OAI211XL U32647 ( .A0(n34458), .A1(n29054), .B0(n34408), .C0(n29053), .Y(
        n15224) );
  XOR2XL U32648 ( .A(n29056), .B(n29055), .Y(n29058) );
  NAND2XL U32649 ( .A(conv_2[394]), .B(n29058), .Y(n29057) );
  OAI211XL U32650 ( .A0(conv_2[394]), .A1(n29058), .B0(n34028), .C0(n29057), 
        .Y(n29059) );
  OAI211XL U32651 ( .A0(n36031), .A1(n29060), .B0(n34408), .C0(n29059), .Y(
        n15213) );
  INVXL U32652 ( .A(conv_2[274]), .Y(n29067) );
  AOI21XL U32653 ( .A0(n29063), .A1(n29062), .B0(n29061), .Y(n29065) );
  NAND2XL U32654 ( .A(conv_2[274]), .B(n29065), .Y(n29064) );
  OAI211XL U32655 ( .A0(conv_2[274]), .A1(n29065), .B0(n36020), .C0(n29064), 
        .Y(n29066) );
  OAI211XL U32656 ( .A0(n30994), .A1(n29067), .B0(n34408), .C0(n29066), .Y(
        n15221) );
  NOR2X1 U32657 ( .A(n29070), .B(n29071), .Y(n31561) );
  AOI21XL U32658 ( .A0(n29071), .A1(n29070), .B0(n31561), .Y(n29072) );
  OAI21XL U32659 ( .A0(n16655), .A1(n29072), .B0(n35630), .Y(n29073) );
  AOI22XL U32660 ( .A0(n33788), .A1(n31560), .B0(conv_3[169]), .B1(n29073), 
        .Y(n29074) );
  NAND2XL U32661 ( .A(n29074), .B(n34097), .Y(n15768) );
  NAND2XL U32662 ( .A(n29076), .B(n29075), .Y(n29078) );
  NAND2XL U32663 ( .A(n29080), .B(n29078), .Y(n29077) );
  OAI211XL U32664 ( .A0(n29080), .A1(n29078), .B0(n33778), .C0(n29077), .Y(
        n29079) );
  OAI211XL U32665 ( .A0(n30412), .A1(n29080), .B0(n34669), .C0(n29079), .Y(
        n15193) );
  OAI2BB1XL U32666 ( .A0N(n33620), .A1N(n29082), .B0(n29081), .Y(n29084) );
  NAND2XL U32667 ( .A(n29086), .B(n29084), .Y(n29083) );
  OAI211XL U32668 ( .A0(n29086), .A1(n29084), .B0(n33982), .C0(n29083), .Y(
        n29085) );
  OAI211XL U32669 ( .A0(n30412), .A1(n29086), .B0(n33815), .C0(n29085), .Y(
        n15192) );
  AOI21XL U32670 ( .A0(n29095), .A1(n29088), .B0(n29087), .Y(n29090) );
  NAND2XL U32671 ( .A(conv_2[532]), .B(n29090), .Y(n29089) );
  OAI211XL U32672 ( .A0(conv_2[532]), .A1(n29090), .B0(n32052), .C0(n29089), 
        .Y(n29091) );
  OAI211XL U32673 ( .A0(n34496), .A1(n29092), .B0(n35859), .C0(n29091), .Y(
        n14851) );
  AOI21XL U32674 ( .A0(n29095), .A1(n29094), .B0(n29093), .Y(n29097) );
  NAND2XL U32675 ( .A(conv_2[534]), .B(n29097), .Y(n29096) );
  OAI211XL U32676 ( .A0(conv_2[534]), .A1(n29097), .B0(n32611), .C0(n29096), 
        .Y(n29098) );
  OAI211XL U32677 ( .A0(n34496), .A1(n29099), .B0(n34735), .C0(n29098), .Y(
        n14849) );
  INVXL U32678 ( .A(conv_2[536]), .Y(n29105) );
  NAND2XL U32679 ( .A(conv_2[536]), .B(n29103), .Y(n29102) );
  OAI211XL U32680 ( .A0(conv_2[536]), .A1(n29103), .B0(n33712), .C0(n29102), 
        .Y(n29104) );
  OAI211XL U32681 ( .A0(n34496), .A1(n29105), .B0(n33815), .C0(n29104), .Y(
        n14847) );
  AOI2BB1XL U32682 ( .A0N(n33480), .A1N(n29107), .B0(n29106), .Y(n29109) );
  NAND2XL U32683 ( .A(conv_3[262]), .B(n29109), .Y(n29108) );
  OAI211XL U32684 ( .A0(conv_3[262]), .A1(n29109), .B0(n36020), .C0(n29108), 
        .Y(n29110) );
  OAI211XL U32685 ( .A0(n35713), .A1(n29111), .B0(n16649), .C0(n29110), .Y(
        n15571) );
  NOR2BXL U32686 ( .AN(n29113), .B(n29112), .Y(n29115) );
  NAND2XL U32687 ( .A(conv_3[260]), .B(n29115), .Y(n29114) );
  OAI211XL U32688 ( .A0(conv_3[260]), .A1(n29115), .B0(n36020), .C0(n29114), 
        .Y(n29116) );
  OAI211XL U32689 ( .A0(n35713), .A1(n29117), .B0(n16649), .C0(n29116), .Y(
        n15573) );
  OAI2BB1XL U32690 ( .A0N(conv_3[250]), .A1N(n29118), .B0(n35700), .Y(n35708)
         );
  NAND4XL U32691 ( .A(conv_3[251]), .B(conv_3[252]), .C(n35700), .D(n35708), 
        .Y(n29125) );
  NAND3XL U32692 ( .A(n35709), .B(n35693), .C(n29182), .Y(n29124) );
  NAND2XL U32693 ( .A(n29125), .B(n29124), .Y(n29121) );
  NAND2XL U32694 ( .A(conv_3[253]), .B(n29121), .Y(n29120) );
  OAI211XL U32695 ( .A0(conv_3[253]), .A1(n29121), .B0(n24378), .C0(n29120), 
        .Y(n29122) );
  OAI211XL U32696 ( .A0(n35706), .A1(n29123), .B0(n35588), .C0(n29122), .Y(
        n15575) );
  AOI22XL U32697 ( .A0(conv_3[253]), .A1(n29125), .B0(n29124), .B1(n29123), 
        .Y(n29127) );
  NAND2XL U32698 ( .A(conv_3[254]), .B(n29127), .Y(n29126) );
  OAI211XL U32699 ( .A0(conv_3[254]), .A1(n29127), .B0(n33982), .C0(n29126), 
        .Y(n29128) );
  OAI211XL U32700 ( .A0(n34676), .A1(n29129), .B0(n35588), .C0(n29128), .Y(
        n15574) );
  AOI21XL U32701 ( .A0(n33478), .A1(n29131), .B0(n29130), .Y(n29133) );
  NAND2XL U32702 ( .A(conv_3[261]), .B(n29133), .Y(n29132) );
  OAI211XL U32703 ( .A0(conv_3[261]), .A1(n29133), .B0(n31735), .C0(n29132), 
        .Y(n29134) );
  OAI211XL U32704 ( .A0(n35713), .A1(n29135), .B0(n16649), .C0(n29134), .Y(
        n15572) );
  OAI21XL U32705 ( .A0(conv_2[229]), .A1(n29138), .B0(n29137), .Y(n29139) );
  AND2XL U32706 ( .A(n33096), .B(n29139), .Y(n29513) );
  AOI2BB1XL U32707 ( .A0N(n29517), .A1N(n29513), .B0(n32876), .Y(n29174) );
  NAND2XL U32708 ( .A(conv_2[233]), .B(n29184), .Y(n29155) );
  OAI31XL U32709 ( .A0(conv_2[233]), .A1(n29184), .A2(conv_2[234]), .B0(n32876), .Y(n29596) );
  OAI21XL U32710 ( .A0(n32876), .A1(n29598), .B0(n29596), .Y(n29141) );
  NAND2XL U32711 ( .A(n29597), .B(n29141), .Y(n29140) );
  OAI211XL U32712 ( .A0(n29597), .A1(n29141), .B0(n16657), .C0(n29140), .Y(
        n29142) );
  OAI211XL U32713 ( .A0(n34458), .A1(n29597), .B0(n34669), .C0(n29142), .Y(
        n15048) );
  AOI21XL U32714 ( .A0(n29455), .A1(n29144), .B0(n29143), .Y(n29146) );
  NAND2XL U32715 ( .A(conv_2[246]), .B(n29146), .Y(n29145) );
  OAI211XL U32716 ( .A0(conv_2[246]), .A1(n29146), .B0(n32660), .C0(n29145), 
        .Y(n29147) );
  OAI211XL U32717 ( .A0(n35945), .A1(n29148), .B0(n33815), .C0(n29147), .Y(
        n15042) );
  AOI21XL U32718 ( .A0(n29455), .A1(n29150), .B0(n29149), .Y(n29152) );
  NAND2XL U32719 ( .A(conv_2[248]), .B(n29152), .Y(n29151) );
  OAI211XL U32720 ( .A0(conv_2[248]), .A1(n29152), .B0(n33778), .C0(n29151), 
        .Y(n29153) );
  OAI211XL U32721 ( .A0(n35945), .A1(n29154), .B0(n34735), .C0(n29153), .Y(
        n15040) );
  OAI32XL U32722 ( .A0(n33096), .A1(n29184), .A2(conv_2[233]), .B0(n32876), 
        .B1(n29155), .Y(n29157) );
  NAND2XL U32723 ( .A(conv_2[234]), .B(n29157), .Y(n29156) );
  OAI211XL U32724 ( .A0(conv_2[234]), .A1(n29157), .B0(n30090), .C0(n29156), 
        .Y(n29158) );
  OAI211XL U32725 ( .A0(n34458), .A1(n29159), .B0(n34735), .C0(n29158), .Y(
        n15049) );
  INVXL U32726 ( .A(conv_3[232]), .Y(n32099) );
  NAND2XL U32727 ( .A(conv_3[231]), .B(n32089), .Y(n32095) );
  NAND2XL U32728 ( .A(conv_3[233]), .B(n35672), .Y(n30690) );
  AOI2BB1XL U32729 ( .A0N(n35673), .A1N(n31061), .B0(n31060), .Y(n29164) );
  NAND2XL U32730 ( .A(conv_3[235]), .B(n29164), .Y(n29163) );
  OAI211XL U32731 ( .A0(conv_3[235]), .A1(n29164), .B0(n32611), .C0(n29163), 
        .Y(n29165) );
  OAI211XL U32732 ( .A0(n35676), .A1(n29166), .B0(n33468), .C0(n29165), .Y(
        n15588) );
  INVXL U32733 ( .A(conv_2[247]), .Y(n29172) );
  AOI2BB1XL U32734 ( .A0N(n35942), .A1N(n29168), .B0(n29167), .Y(n29170) );
  NAND2XL U32735 ( .A(conv_2[247]), .B(n29170), .Y(n29169) );
  OAI211XL U32736 ( .A0(conv_2[247]), .A1(n29170), .B0(n34028), .C0(n29169), 
        .Y(n29171) );
  OAI211XL U32737 ( .A0(n35945), .A1(n29172), .B0(n33815), .C0(n29171), .Y(
        n15041) );
  NAND2XL U32738 ( .A(conv_2[231]), .B(n29176), .Y(n29175) );
  OAI211XL U32739 ( .A0(conv_2[231]), .A1(n29176), .B0(n27932), .C0(n29175), 
        .Y(n29177) );
  OAI211XL U32740 ( .A0(n34458), .A1(n29178), .B0(n35859), .C0(n29177), .Y(
        n15052) );
  AOI32XL U32741 ( .A0(conv_3[251]), .A1(n35700), .A2(n35708), .B0(n35693), 
        .B1(n35709), .Y(n29180) );
  NAND2XL U32742 ( .A(n29182), .B(n29180), .Y(n29179) );
  OAI211XL U32743 ( .A0(n29182), .A1(n29180), .B0(n33778), .C0(n29179), .Y(
        n29181) );
  OAI211XL U32744 ( .A0(n35706), .A1(n29182), .B0(n33468), .C0(n29181), .Y(
        n15576) );
  AOI21XL U32745 ( .A0(n29184), .A1(n32876), .B0(n29183), .Y(n29186) );
  NAND2XL U32746 ( .A(conv_2[233]), .B(n29186), .Y(n29185) );
  OAI211XL U32747 ( .A0(conv_2[233]), .A1(n29186), .B0(n33982), .C0(n29185), 
        .Y(n29187) );
  OAI211XL U32748 ( .A0(n34458), .A1(n29188), .B0(n33815), .C0(n29187), .Y(
        n15050) );
  INVXL U32749 ( .A(conv_1[535]), .Y(n29194) );
  NAND2XL U32750 ( .A(conv_1[535]), .B(n29192), .Y(n29191) );
  OAI211XL U32751 ( .A0(conv_1[535]), .A1(n29192), .B0(n33778), .C0(n29191), 
        .Y(n29193) );
  OAI211XL U32752 ( .A0(n33432), .A1(n29194), .B0(n34689), .C0(n29193), .Y(
        n15928) );
  AOI21XL U32753 ( .A0(n29281), .A1(conv_1[263]), .B0(n30191), .Y(n29227) );
  NAND2XL U32754 ( .A(conv_1[264]), .B(n29199), .Y(n29198) );
  OAI211XL U32755 ( .A0(conv_1[264]), .A1(n29199), .B0(n33778), .C0(n29198), 
        .Y(n29200) );
  OAI211XL U32756 ( .A0(n34080), .A1(n29201), .B0(n34544), .C0(n29200), .Y(
        n16199) );
  AOI2BB1XL U32757 ( .A0N(n30191), .A1N(n29203), .B0(n29202), .Y(n29205) );
  NAND2XL U32758 ( .A(conv_1[261]), .B(n29205), .Y(n29204) );
  OAI211XL U32759 ( .A0(conv_1[261]), .A1(n29205), .B0(n34028), .C0(n29204), 
        .Y(n29206) );
  OAI211XL U32760 ( .A0(n34080), .A1(n29207), .B0(n16652), .C0(n29206), .Y(
        n16202) );
  OAI2BB1XL U32761 ( .A0N(n29216), .A1N(n29209), .B0(n29208), .Y(n29211) );
  NAND2XL U32762 ( .A(n29213), .B(n29211), .Y(n29210) );
  OAI211XL U32763 ( .A0(n29213), .A1(n29211), .B0(n33778), .C0(n29210), .Y(
        n29212) );
  OAI211XL U32764 ( .A0(n33432), .A1(n29213), .B0(n16652), .C0(n29212), .Y(
        n15931) );
  AOI2BB1XL U32765 ( .A0N(n29216), .A1N(n29215), .B0(n29214), .Y(n29218) );
  NAND2XL U32766 ( .A(conv_1[534]), .B(n29218), .Y(n29217) );
  OAI211XL U32767 ( .A0(conv_1[534]), .A1(n29218), .B0(n31735), .C0(n29217), 
        .Y(n29219) );
  OAI211XL U32768 ( .A0(n33432), .A1(n29220), .B0(n34682), .C0(n29219), .Y(
        n15929) );
  INVXL U32769 ( .A(conv_1[432]), .Y(n29329) );
  OAI2BB1XL U32770 ( .A0N(conv_1[431]), .A1N(n35508), .B0(n29328), .Y(n29327)
         );
  OAI21XL U32771 ( .A0(n29330), .A1(n29328), .B0(n29327), .Y(n29225) );
  NAND2XL U32772 ( .A(n29329), .B(n29225), .Y(n29224) );
  OAI211XL U32773 ( .A0(n29329), .A1(n29225), .B0(n16656), .C0(n29224), .Y(
        n29226) );
  OAI211XL U32774 ( .A0(n35504), .A1(n29329), .B0(n34696), .C0(n29226), .Y(
        n16031) );
  NAND4XL U32775 ( .A(conv_1[266]), .B(conv_1[267]), .C(n29350), .D(n29229), 
        .Y(n34079) );
  NAND4BXL U32776 ( .AN(n29350), .B(n30191), .C(n29355), .D(n29326), .Y(n34078) );
  AOI22XL U32777 ( .A0(conv_1[268]), .A1(n34079), .B0(n34078), .B1(n34083), 
        .Y(n29231) );
  NAND2XL U32778 ( .A(conv_1[269]), .B(n29231), .Y(n29230) );
  OAI211XL U32779 ( .A0(conv_1[269]), .A1(n29231), .B0(n16657), .C0(n29230), 
        .Y(n29232) );
  OAI211XL U32780 ( .A0(n33442), .A1(n29233), .B0(n16652), .C0(n29232), .Y(
        n16194) );
  AOI21XL U32781 ( .A0(n29236), .A1(n29235), .B0(n29234), .Y(n29238) );
  NAND2XL U32782 ( .A(conv_1[533]), .B(n29238), .Y(n29237) );
  OAI211XL U32783 ( .A0(conv_1[533]), .A1(n29238), .B0(n24378), .C0(n29237), 
        .Y(n29239) );
  OAI211XL U32784 ( .A0(n33432), .A1(n29240), .B0(n34544), .C0(n29239), .Y(
        n15930) );
  OAI211XL U32785 ( .A0(n29242), .A1(conv_1[531]), .B0(n33822), .C0(n29241), 
        .Y(n29243) );
  OAI211XL U32786 ( .A0(n33432), .A1(n29244), .B0(n34682), .C0(n29243), .Y(
        n15932) );
  NAND4XL U32787 ( .A(conv_1[521]), .B(conv_1[522]), .C(n30267), .D(n35550), 
        .Y(n30257) );
  NAND3XL U32788 ( .A(n35551), .B(n29246), .C(n29245), .Y(n30256) );
  AOI22XL U32789 ( .A0(conv_1[523]), .A1(n30257), .B0(n30256), .B1(n30261), 
        .Y(n29248) );
  NAND2XL U32790 ( .A(conv_1[524]), .B(n29248), .Y(n29247) );
  OAI211XL U32791 ( .A0(conv_1[524]), .A1(n29248), .B0(n33778), .C0(n29247), 
        .Y(n29249) );
  OAI211XL U32792 ( .A0(n33853), .A1(n29250), .B0(n34689), .C0(n29249), .Y(
        n15939) );
  AOI22XL U32793 ( .A0(conv_1[283]), .A1(n29253), .B0(n29252), .B1(n29251), 
        .Y(n29255) );
  NAND2XL U32794 ( .A(conv_1[284]), .B(n29255), .Y(n29254) );
  OAI211XL U32795 ( .A0(conv_1[284]), .A1(n29255), .B0(n33712), .C0(n29254), 
        .Y(n29256) );
  OAI211XL U32796 ( .A0(n33442), .A1(n29257), .B0(n34682), .C0(n29256), .Y(
        n16179) );
  NAND2XL U32797 ( .A(conv_1[113]), .B(n31343), .Y(n31342) );
  NAND4XL U32798 ( .A(conv_1[116]), .B(conv_1[117]), .C(n31344), .D(n35332), 
        .Y(n33239) );
  OAI31XL U32799 ( .A0(conv_1[113]), .A1(conv_1[114]), .A2(n31343), .B0(n34557), .Y(n34555) );
  OAI2BB1XL U32800 ( .A0N(n34561), .A1N(n34555), .B0(n34557), .Y(n35331) );
  NAND3XL U32801 ( .A(n35333), .B(n34557), .C(n29338), .Y(n33238) );
  INVXL U32802 ( .A(conv_1[118]), .Y(n33242) );
  AOI22XL U32803 ( .A0(conv_1[118]), .A1(n33239), .B0(n33238), .B1(n33242), 
        .Y(n29259) );
  NAND2XL U32804 ( .A(conv_1[119]), .B(n29259), .Y(n29258) );
  OAI211XL U32805 ( .A0(conv_1[119]), .A1(n29259), .B0(n32181), .C0(n29258), 
        .Y(n29260) );
  OAI211XL U32806 ( .A0(n34676), .A1(n29261), .B0(n34281), .C0(n29260), .Y(
        n16344) );
  AOI2BB1XL U32807 ( .A0N(n35404), .A1N(n29263), .B0(n29262), .Y(n29265) );
  NAND2XL U32808 ( .A(conv_1[231]), .B(n29265), .Y(n29264) );
  OAI211XL U32809 ( .A0(conv_1[231]), .A1(n29265), .B0(n27932), .C0(n29264), 
        .Y(n29266) );
  OAI211XL U32810 ( .A0(n35408), .A1(n29267), .B0(n16652), .C0(n29266), .Y(
        n16232) );
  AOI2BB1XL U32811 ( .A0N(n33654), .A1N(n29269), .B0(n29268), .Y(n29271) );
  NAND2XL U32812 ( .A(conv_1[396]), .B(n29271), .Y(n29270) );
  OAI211XL U32813 ( .A0(conv_1[396]), .A1(n29271), .B0(n33822), .C0(n29270), 
        .Y(n29272) );
  OAI211XL U32814 ( .A0(n35477), .A1(n29273), .B0(n34281), .C0(n29272), .Y(
        n16067) );
  NAND2XL U32815 ( .A(conv_1[395]), .B(n29277), .Y(n29276) );
  OAI211XL U32816 ( .A0(conv_1[395]), .A1(n29277), .B0(n33822), .C0(n29276), 
        .Y(n29278) );
  OAI211XL U32817 ( .A0(n35477), .A1(n29279), .B0(n16652), .C0(n29278), .Y(
        n16068) );
  INVXL U32818 ( .A(conv_1[263]), .Y(n29285) );
  AOI2BB1XL U32819 ( .A0N(n30191), .A1N(n29281), .B0(n29280), .Y(n29283) );
  NAND2XL U32820 ( .A(conv_1[263]), .B(n29283), .Y(n29282) );
  OAI211XL U32821 ( .A0(conv_1[263]), .A1(n29283), .B0(n34666), .C0(n29282), 
        .Y(n29284) );
  OAI211XL U32822 ( .A0(n34080), .A1(n29285), .B0(n34696), .C0(n29284), .Y(
        n16200) );
  AOI21XL U32823 ( .A0(n34775), .A1(n29287), .B0(n29286), .Y(n29289) );
  NAND2XL U32824 ( .A(conv_1[411]), .B(n29289), .Y(n29288) );
  OAI211XL U32825 ( .A0(conv_1[411]), .A1(n29289), .B0(n34028), .C0(n29288), 
        .Y(n29290) );
  OAI211XL U32826 ( .A0(n35487), .A1(n29291), .B0(n34696), .C0(n29290), .Y(
        n16052) );
  NAND2XL U32827 ( .A(conv_1[110]), .B(n29295), .Y(n29294) );
  OAI211XL U32828 ( .A0(conv_1[110]), .A1(n29295), .B0(n32181), .C0(n29294), 
        .Y(n29296) );
  OAI211XL U32829 ( .A0(n35330), .A1(n29297), .B0(n34696), .C0(n29296), .Y(
        n16353) );
  NAND2XL U32830 ( .A(conv_1[415]), .B(n29301), .Y(n29300) );
  OAI211XL U32831 ( .A0(conv_1[415]), .A1(n29301), .B0(n32181), .C0(n29300), 
        .Y(n29302) );
  OAI211XL U32832 ( .A0(n35487), .A1(n29303), .B0(n34281), .C0(n29302), .Y(
        n16048) );
  INVXL U32833 ( .A(conv_1[125]), .Y(n29309) );
  NAND2XL U32834 ( .A(conv_1[125]), .B(n29307), .Y(n29306) );
  OAI211XL U32835 ( .A0(conv_1[125]), .A1(n29307), .B0(n32181), .C0(n29306), 
        .Y(n29308) );
  OAI211XL U32836 ( .A0(n34296), .A1(n29309), .B0(n34682), .C0(n29308), .Y(
        n16338) );
  NAND2XL U32837 ( .A(conv_1[290]), .B(n29313), .Y(n29312) );
  OAI211XL U32838 ( .A0(conv_1[290]), .A1(n29313), .B0(n34028), .C0(n29312), 
        .Y(n29314) );
  OAI211XL U32839 ( .A0(n34325), .A1(n29315), .B0(n34281), .C0(n29314), .Y(
        n16173) );
  AOI21XL U32840 ( .A0(n29339), .A1(n29317), .B0(n29316), .Y(n29319) );
  NAND2XL U32841 ( .A(conv_1[276]), .B(n29319), .Y(n29318) );
  OAI211XL U32842 ( .A0(conv_1[276]), .A1(n29319), .B0(n16656), .C0(n29318), 
        .Y(n29320) );
  OAI211XL U32843 ( .A0(n35426), .A1(n29321), .B0(n34544), .C0(n29320), .Y(
        n16187) );
  AOI21XL U32844 ( .A0(n29350), .A1(n30191), .B0(n29322), .Y(n29324) );
  NAND2XL U32845 ( .A(conv_1[266]), .B(n29324), .Y(n29323) );
  OAI211XL U32846 ( .A0(conv_1[266]), .A1(n29324), .B0(n32656), .C0(n29323), 
        .Y(n29325) );
  OAI211XL U32847 ( .A0(n34080), .A1(n29326), .B0(n16652), .C0(n29325), .Y(
        n16197) );
  NAND3XL U32848 ( .A(conv_1[432]), .B(n29328), .C(n29327), .Y(n29396) );
  NAND3XL U32849 ( .A(intadd_1_B_2_), .B(n29330), .C(n29329), .Y(n29395) );
  INVXL U32850 ( .A(conv_1[433]), .Y(n29400) );
  AOI22XL U32851 ( .A0(conv_1[433]), .A1(n29396), .B0(n29395), .B1(n29400), 
        .Y(n29332) );
  NAND2XL U32852 ( .A(conv_1[434]), .B(n29332), .Y(n29331) );
  OAI211XL U32853 ( .A0(conv_1[434]), .A1(n29332), .B0(n28751), .C0(n29331), 
        .Y(n29333) );
  OAI211XL U32854 ( .A0(n33853), .A1(n29334), .B0(n34544), .C0(n29333), .Y(
        n16029) );
  AOI32XL U32855 ( .A0(conv_1[116]), .A1(n31344), .A2(n35332), .B0(n34557), 
        .B1(n35333), .Y(n29336) );
  NAND2XL U32856 ( .A(n29338), .B(n29336), .Y(n29335) );
  OAI211XL U32857 ( .A0(n29338), .A1(n29336), .B0(n32181), .C0(n29335), .Y(
        n29337) );
  OAI211XL U32858 ( .A0(n35330), .A1(n29338), .B0(n16652), .C0(n29337), .Y(
        n16346) );
  AOI32XL U32859 ( .A0(conv_1[281]), .A1(n29339), .A2(n35428), .B0(n29364), 
        .B1(n35429), .Y(n29341) );
  NAND2XL U32860 ( .A(n29343), .B(n29341), .Y(n29340) );
  OAI211XL U32861 ( .A0(n29343), .A1(n29341), .B0(n16656), .C0(n29340), .Y(
        n29342) );
  OAI211XL U32862 ( .A0(n35426), .A1(n29343), .B0(n34281), .C0(n29342), .Y(
        n16181) );
  INVXL U32863 ( .A(conv_1[277]), .Y(n29349) );
  AOI2BB1XL U32864 ( .A0N(n29364), .A1N(n29345), .B0(n29344), .Y(n29347) );
  NAND2XL U32865 ( .A(conv_1[277]), .B(n29347), .Y(n29346) );
  OAI211XL U32866 ( .A0(conv_1[277]), .A1(n29347), .B0(n31735), .C0(n29346), 
        .Y(n29348) );
  OAI211XL U32867 ( .A0(n35426), .A1(n29349), .B0(n34696), .C0(n29348), .Y(
        n16186) );
  OAI21XL U32868 ( .A0(conv_1[266]), .A1(n29350), .B0(n30191), .Y(n29351) );
  AOI32XL U32869 ( .A0(conv_1[266]), .A1(n29351), .A2(n29350), .B0(n30191), 
        .B1(n29351), .Y(n29353) );
  NAND2XL U32870 ( .A(n29355), .B(n29353), .Y(n29352) );
  OAI211XL U32871 ( .A0(n29355), .A1(n29353), .B0(n32611), .C0(n29352), .Y(
        n29354) );
  OAI211XL U32872 ( .A0(n34080), .A1(n29355), .B0(n34696), .C0(n29354), .Y(
        n16196) );
  AOI2BB1XL U32873 ( .A0N(n33654), .A1N(n31279), .B0(n31280), .Y(n29360) );
  NAND2XL U32874 ( .A(conv_1[398]), .B(n29360), .Y(n29359) );
  OAI211XL U32875 ( .A0(conv_1[398]), .A1(n29360), .B0(n33822), .C0(n29359), 
        .Y(n29361) );
  OAI211XL U32876 ( .A0(n35477), .A1(n29362), .B0(n16652), .C0(n29361), .Y(
        n16065) );
  INVXL U32877 ( .A(conv_1[280]), .Y(n29369) );
  AOI21XL U32878 ( .A0(n29365), .A1(n29364), .B0(n29363), .Y(n29367) );
  NAND2XL U32879 ( .A(conv_1[280]), .B(n29367), .Y(n29366) );
  OAI211XL U32880 ( .A0(conv_1[280]), .A1(n29367), .B0(n24499), .C0(n29366), 
        .Y(n29368) );
  OAI211XL U32881 ( .A0(n35426), .A1(n29369), .B0(n16652), .C0(n29368), .Y(
        n16183) );
  INVXL U32882 ( .A(conv_1[275]), .Y(n29375) );
  NOR2BXL U32883 ( .AN(n29371), .B(n29370), .Y(n29373) );
  NAND2XL U32884 ( .A(conv_1[275]), .B(n29373), .Y(n29372) );
  OAI211XL U32885 ( .A0(conv_1[275]), .A1(n29373), .B0(n33712), .C0(n29372), 
        .Y(n29374) );
  OAI211XL U32886 ( .A0(n35426), .A1(n29375), .B0(n34689), .C0(n29374), .Y(
        n16188) );
  INVXL U32887 ( .A(conv_1[291]), .Y(n29381) );
  AOI2BB1XL U32888 ( .A0N(n34319), .A1N(n29377), .B0(n29376), .Y(n29379) );
  NAND2XL U32889 ( .A(conv_1[291]), .B(n29379), .Y(n29378) );
  OAI211XL U32890 ( .A0(conv_1[291]), .A1(n29379), .B0(n33712), .C0(n29378), 
        .Y(n29380) );
  OAI211XL U32891 ( .A0(n34325), .A1(n29381), .B0(n16652), .C0(n29380), .Y(
        n16172) );
  INVXL U32892 ( .A(conv_1[321]), .Y(n29389) );
  AOI2BB1XL U32893 ( .A0N(n29383), .A1N(conv_1[320]), .B0(n29382), .Y(n29384)
         );
  AOI2BB1XL U32894 ( .A0N(n34259), .A1N(n29385), .B0(n29384), .Y(n29387) );
  NAND2XL U32895 ( .A(conv_1[321]), .B(n29387), .Y(n29386) );
  OAI211XL U32896 ( .A0(conv_1[321]), .A1(n29387), .B0(n32660), .C0(n29386), 
        .Y(n29388) );
  OAI211XL U32897 ( .A0(n34263), .A1(n29389), .B0(n34689), .C0(n29388), .Y(
        n16142) );
  AOI21XL U32898 ( .A0(n34289), .A1(n34292), .B0(n29390), .Y(n29392) );
  NAND2XL U32899 ( .A(conv_1[127]), .B(n29392), .Y(n29391) );
  OAI211XL U32900 ( .A0(conv_1[127]), .A1(n29392), .B0(n32181), .C0(n29391), 
        .Y(n29393) );
  OAI211XL U32901 ( .A0(n34296), .A1(n29394), .B0(n34689), .C0(n29393), .Y(
        n16336) );
  NAND2XL U32902 ( .A(n29396), .B(n29395), .Y(n29398) );
  NAND2XL U32903 ( .A(conv_1[433]), .B(n29398), .Y(n29397) );
  OAI211XL U32904 ( .A0(conv_1[433]), .A1(n29398), .B0(n28751), .C0(n29397), 
        .Y(n29399) );
  OAI211XL U32905 ( .A0(n35504), .A1(n29400), .B0(n34682), .C0(n29399), .Y(
        n16030) );
  INVXL U32906 ( .A(conv_1[427]), .Y(n29406) );
  AOI2BB1XL U32907 ( .A0N(intadd_1_B_2_), .A1N(n29402), .B0(n29401), .Y(n29404) );
  NAND2XL U32908 ( .A(conv_1[427]), .B(n29404), .Y(n29403) );
  OAI211XL U32909 ( .A0(conv_1[427]), .A1(n29404), .B0(n32181), .C0(n29403), 
        .Y(n29405) );
  OAI211XL U32910 ( .A0(n35504), .A1(n29406), .B0(n34696), .C0(n29405), .Y(
        n16036) );
  AOI21XL U32911 ( .A0(n29409), .A1(n29408), .B0(n29407), .Y(n29411) );
  NAND2XL U32912 ( .A(conv_2[259]), .B(n29411), .Y(n29410) );
  OAI211XL U32913 ( .A0(conv_2[259]), .A1(n29411), .B0(n32181), .C0(n29410), 
        .Y(n29412) );
  OAI211XL U32914 ( .A0(n34601), .A1(n29413), .B0(n34408), .C0(n29412), .Y(
        n15222) );
  NAND2XL U32915 ( .A(conv_3[258]), .B(n29417), .Y(n29416) );
  OAI211XL U32916 ( .A0(conv_3[258]), .A1(n29417), .B0(n32611), .C0(n29416), 
        .Y(n29418) );
  OAI211XL U32917 ( .A0(n35713), .A1(n29419), .B0(n29418), .C0(n35574), .Y(
        n15798) );
  NOR2BXL U32918 ( .AN(n29421), .B(n29420), .Y(n29423) );
  NAND2XL U32919 ( .A(conv_2[408]), .B(n29423), .Y(n29422) );
  OAI211XL U32920 ( .A0(conv_2[408]), .A1(n29423), .B0(n32660), .C0(n29422), 
        .Y(n29424) );
  OAI211XL U32921 ( .A0(n36047), .A1(n29425), .B0(n29424), .C0(n34105), .Y(
        n15248) );
  INVXL U32922 ( .A(conv_3[19]), .Y(n29436) );
  OAI21XL U32923 ( .A0(n30195), .A1(n18997), .B0(n30549), .Y(n29430) );
  INVXL U32924 ( .A(n29430), .Y(n30550) );
  INVXL U32925 ( .A(conv_3[17]), .Y(n30555) );
  OAI22XL U32926 ( .A0(n18997), .A1(n30549), .B0(n30550), .B1(n30555), .Y(
        n29977) );
  NAND2XL U32927 ( .A(conv_3[19]), .B(n29434), .Y(n29433) );
  OAI211XL U32928 ( .A0(conv_3[19]), .A1(n29434), .B0(n34028), .C0(n29433), 
        .Y(n29435) );
  OAI211XL U32929 ( .A0(n35576), .A1(n29436), .B0(n29435), .C0(n34097), .Y(
        n15778) );
  OAI211XL U32930 ( .A0(conv_2[524]), .A1(n29441), .B0(n33982), .C0(n29440), 
        .Y(n29442) );
  NAND2XL U32931 ( .A(conv_2[380]), .B(n29447), .Y(n29446) );
  OAI211XL U32932 ( .A0(conv_2[380]), .A1(n29447), .B0(n34666), .C0(n29446), 
        .Y(n29448) );
  OAI211XL U32933 ( .A0(n36028), .A1(n29449), .B0(n33815), .C0(n29448), .Y(
        n14953) );
  NAND2XL U32934 ( .A(conv_2[338]), .B(n35996), .Y(n35994) );
  NAND4XL U32935 ( .A(conv_2[341]), .B(conv_2[342]), .C(n35997), .D(n36005), 
        .Y(n34218) );
  OAI31XL U32936 ( .A0(conv_2[338]), .A1(conv_2[339]), .A2(n35996), .B0(n35995), .Y(n29610) );
  OAI2BB1XL U32937 ( .A0N(n29615), .A1N(n29610), .B0(n35995), .Y(n36004) );
  INVXL U32938 ( .A(conv_2[342]), .Y(n29505) );
  NAND3XL U32939 ( .A(n36006), .B(n35995), .C(n29505), .Y(n34217) );
  AOI22XL U32940 ( .A0(conv_2[343]), .A1(n34218), .B0(n34217), .B1(n34221), 
        .Y(n29451) );
  NAND2XL U32941 ( .A(conv_2[344]), .B(n29451), .Y(n29450) );
  OAI211XL U32942 ( .A0(conv_2[344]), .A1(n29451), .B0(n27932), .C0(n29450), 
        .Y(n29452) );
  OAI211XL U32943 ( .A0(n33442), .A1(n29453), .B0(n34735), .C0(n29452), .Y(
        n14974) );
  OAI21XL U32944 ( .A0(n29456), .A1(n29455), .B0(n29454), .Y(n29458) );
  NAND2XL U32945 ( .A(n29460), .B(n29458), .Y(n29457) );
  OAI211XL U32946 ( .A0(n29460), .A1(n29458), .B0(n27932), .C0(n29457), .Y(
        n29459) );
  OAI211XL U32947 ( .A0(n35945), .A1(n29460), .B0(n33815), .C0(n29459), .Y(
        n15036) );
  NAND4XL U32948 ( .A(conv_2[356]), .B(conv_2[357]), .C(n33925), .D(n36012), 
        .Y(n29474) );
  NAND3XL U32949 ( .A(n36013), .B(n29526), .C(n29461), .Y(n29473) );
  AOI22XL U32950 ( .A0(conv_2[358]), .A1(n29474), .B0(n29473), .B1(n29478), 
        .Y(n29463) );
  NAND2XL U32951 ( .A(conv_2[359]), .B(n29463), .Y(n29462) );
  OAI211XL U32952 ( .A0(conv_2[359]), .A1(n29463), .B0(n33778), .C0(n29462), 
        .Y(n29464) );
  OAI211XL U32953 ( .A0(n33853), .A1(n29465), .B0(n34735), .C0(n29464), .Y(
        n14964) );
  AOI22XL U32954 ( .A0(conv_2[373]), .A1(n29468), .B0(n29467), .B1(n29466), 
        .Y(n29470) );
  NAND2XL U32955 ( .A(conv_2[374]), .B(n29470), .Y(n29469) );
  OAI211XL U32956 ( .A0(conv_2[374]), .A1(n29470), .B0(n34028), .C0(n29469), 
        .Y(n29471) );
  OAI211XL U32957 ( .A0(n34520), .A1(n29472), .B0(n34669), .C0(n29471), .Y(
        n14954) );
  NAND2XL U32958 ( .A(n29474), .B(n29473), .Y(n29476) );
  NAND2XL U32959 ( .A(conv_2[358]), .B(n29476), .Y(n29475) );
  OAI211XL U32960 ( .A0(conv_2[358]), .A1(n29476), .B0(n16657), .C0(n29475), 
        .Y(n29477) );
  OAI211XL U32961 ( .A0(n36010), .A1(n29478), .B0(n35859), .C0(n29477), .Y(
        n14965) );
  OAI32XL U32962 ( .A0(n29526), .A1(n29481), .A2(n29480), .B0(n33925), .B1(
        n29479), .Y(n29483) );
  NAND2XL U32963 ( .A(conv_2[355]), .B(n29483), .Y(n29482) );
  OAI211XL U32964 ( .A0(conv_2[355]), .A1(n29483), .B0(n33778), .C0(n29482), 
        .Y(n29484) );
  OAI211XL U32965 ( .A0(n36010), .A1(n29485), .B0(n33815), .C0(n29484), .Y(
        n14968) );
  AOI21XL U32966 ( .A0(n33321), .A1(n29487), .B0(n29486), .Y(n29489) );
  NAND2XL U32967 ( .A(conv_2[411]), .B(n29489), .Y(n29488) );
  OAI211XL U32968 ( .A0(conv_2[411]), .A1(n29489), .B0(n24499), .C0(n29488), 
        .Y(n29490) );
  OAI211XL U32969 ( .A0(n36047), .A1(n29491), .B0(n35859), .C0(n29490), .Y(
        n14932) );
  INVXL U32970 ( .A(conv_2[369]), .Y(n29497) );
  NAND2XL U32971 ( .A(conv_2[369]), .B(n29495), .Y(n29494) );
  OAI211XL U32972 ( .A0(conv_2[369]), .A1(n29495), .B0(n33778), .C0(n29494), 
        .Y(n29496) );
  OAI211XL U32973 ( .A0(n36017), .A1(n29497), .B0(n34735), .C0(n29496), .Y(
        n14959) );
  OAI21XL U32974 ( .A0(conv_2[398]), .A1(n34635), .B0(n34634), .Y(n34636) );
  NAND2XL U32975 ( .A(n34640), .B(n34636), .Y(n33142) );
  AOI31XL U32976 ( .A0(conv_2[399]), .A1(conv_2[398]), .A2(n34635), .B0(n34634), .Y(n33141) );
  AOI21XL U32977 ( .A0(n34634), .A1(n33142), .B0(n33141), .Y(n29500) );
  NAND2XL U32978 ( .A(conv_2[400]), .B(n29500), .Y(n29499) );
  OAI211XL U32979 ( .A0(conv_2[400]), .A1(n29500), .B0(n33712), .C0(n29499), 
        .Y(n29501) );
  OAI211XL U32980 ( .A0(n36031), .A1(n33140), .B0(n33815), .C0(n29501), .Y(
        n14938) );
  AOI32XL U32981 ( .A0(conv_2[341]), .A1(n35997), .A2(n36005), .B0(n35995), 
        .B1(n36006), .Y(n29503) );
  NAND2XL U32982 ( .A(n29505), .B(n29503), .Y(n29502) );
  OAI211XL U32983 ( .A0(n29505), .A1(n29503), .B0(n16657), .C0(n29502), .Y(
        n29504) );
  OAI211XL U32984 ( .A0(n36003), .A1(n29505), .B0(n34735), .C0(n29504), .Y(
        n14976) );
  INVXL U32985 ( .A(conv_2[368]), .Y(n29511) );
  AOI21XL U32986 ( .A0(n29507), .A1(n34570), .B0(n29506), .Y(n29509) );
  NAND2XL U32987 ( .A(conv_2[368]), .B(n29509), .Y(n29508) );
  OAI211XL U32988 ( .A0(conv_2[368]), .A1(n29509), .B0(n33778), .C0(n29508), 
        .Y(n29510) );
  OAI211XL U32989 ( .A0(n36017), .A1(n29511), .B0(n35859), .C0(n29510), .Y(
        n14960) );
  NAND2XL U32990 ( .A(conv_2[230]), .B(n29515), .Y(n29514) );
  OAI211XL U32991 ( .A0(conv_2[230]), .A1(n29515), .B0(n34666), .C0(n29514), 
        .Y(n29516) );
  OAI211XL U32992 ( .A0(n34458), .A1(n29517), .B0(n33815), .C0(n29516), .Y(
        n15053) );
  AOI21XL U32993 ( .A0(n29523), .A1(n29526), .B0(n29518), .Y(n29520) );
  NAND2XL U32994 ( .A(conv_2[352]), .B(n29520), .Y(n29519) );
  OAI211XL U32995 ( .A0(conv_2[352]), .A1(n29520), .B0(n36020), .C0(n29519), 
        .Y(n29521) );
  OAI211XL U32996 ( .A0(n36010), .A1(n29522), .B0(n34669), .C0(n29521), .Y(
        n14971) );
  INVXL U32997 ( .A(conv_2[353]), .Y(n29530) );
  AOI2BB1XL U32998 ( .A0N(conv_2[352]), .A1N(n29523), .B0(n33925), .Y(n29524)
         );
  AOI2BB1XL U32999 ( .A0N(n29526), .A1N(n29525), .B0(n29524), .Y(n29528) );
  NAND2XL U33000 ( .A(conv_2[353]), .B(n29528), .Y(n29527) );
  OAI211XL U33001 ( .A0(conv_2[353]), .A1(n29528), .B0(n33982), .C0(n29527), 
        .Y(n29529) );
  OAI211XL U33002 ( .A0(n36010), .A1(n29530), .B0(n35859), .C0(n29529), .Y(
        n14970) );
  INVXL U33003 ( .A(conv_2[398]), .Y(n29535) );
  AOI21XL U33004 ( .A0(n34635), .A1(n34634), .B0(n29531), .Y(n29533) );
  NAND2XL U33005 ( .A(conv_2[398]), .B(n29533), .Y(n29532) );
  OAI211XL U33006 ( .A0(conv_2[398]), .A1(n29533), .B0(n24499), .C0(n29532), 
        .Y(n29534) );
  OAI211XL U33007 ( .A0(n36031), .A1(n29535), .B0(n35859), .C0(n29534), .Y(
        n14940) );
  INVXL U33008 ( .A(conv_2[371]), .Y(n29540) );
  AOI21XL U33009 ( .A0(n34571), .A1(n34570), .B0(n29536), .Y(n29538) );
  NAND2XL U33010 ( .A(conv_2[371]), .B(n29538), .Y(n29537) );
  OAI211XL U33011 ( .A0(conv_2[371]), .A1(n29538), .B0(n24499), .C0(n29537), 
        .Y(n29539) );
  OAI211XL U33012 ( .A0(n36017), .A1(n29540), .B0(n33815), .C0(n29539), .Y(
        n14957) );
  NAND2XL U33013 ( .A(conv_1[498]), .B(n29544), .Y(n29543) );
  OAI211XL U33014 ( .A0(conv_1[498]), .A1(n29544), .B0(n27932), .C0(n29543), 
        .Y(n29545) );
  OAI211XL U33015 ( .A0(n33427), .A1(n29546), .B0(n32867), .C0(n29545), .Y(
        n15965) );
  INVXL U33016 ( .A(conv_2[483]), .Y(n29552) );
  NAND2XL U33017 ( .A(conv_2[483]), .B(n29550), .Y(n29549) );
  OAI211XL U33018 ( .A0(conv_2[483]), .A1(n29550), .B0(n33982), .C0(n29549), 
        .Y(n29551) );
  OAI211XL U33019 ( .A0(n34137), .A1(n29552), .B0(n34105), .C0(n29551), .Y(
        n15243) );
  NAND2XL U33020 ( .A(conv_2[438]), .B(n29556), .Y(n29555) );
  OAI211XL U33021 ( .A0(conv_2[438]), .A1(n29556), .B0(n32660), .C0(n29555), 
        .Y(n29557) );
  OAI211XL U33022 ( .A0(n36070), .A1(n29558), .B0(n34105), .C0(n29557), .Y(
        n15246) );
  INVXL U33023 ( .A(conv_2[468]), .Y(n29564) );
  NOR2BXL U33024 ( .AN(n29560), .B(n29559), .Y(n29562) );
  NAND2XL U33025 ( .A(conv_2[468]), .B(n29562), .Y(n29561) );
  OAI211XL U33026 ( .A0(conv_2[468]), .A1(n29562), .B0(n36020), .C0(n29561), 
        .Y(n29563) );
  OAI211XL U33027 ( .A0(n34177), .A1(n29564), .B0(n34105), .C0(n29563), .Y(
        n15244) );
  NAND2XL U33028 ( .A(conv_2[393]), .B(n29568), .Y(n29567) );
  OAI211XL U33029 ( .A0(conv_2[393]), .A1(n29568), .B0(n32660), .C0(n29567), 
        .Y(n29569) );
  OAI211XL U33030 ( .A0(n36031), .A1(n29570), .B0(n34105), .C0(n29569), .Y(
        n15249) );
  INVXL U33031 ( .A(conv_1[408]), .Y(n29576) );
  NAND2XL U33032 ( .A(conv_1[408]), .B(n29574), .Y(n29573) );
  OAI211XL U33033 ( .A0(conv_1[408]), .A1(n29574), .B0(n32181), .C0(n29573), 
        .Y(n29575) );
  OAI211XL U33034 ( .A0(n35487), .A1(n29576), .B0(n32867), .C0(n29575), .Y(
        n16055) );
  AOI22XL U33035 ( .A0(n30090), .A1(n29579), .B0(conv_2[491]), .B1(n33598), 
        .Y(n29580) );
  NAND2XL U33036 ( .A(n29580), .B(n35859), .Y(n14877) );
  OAI2BB1XL U33037 ( .A0N(n29583), .A1N(n29582), .B0(n29581), .Y(n29585) );
  AOI211XL U33038 ( .A0(n29587), .A1(n29585), .B0(n36001), .C0(n29584), .Y(
        n29586) );
  AOI2BB1XL U33039 ( .A0N(n29587), .A1N(n30958), .B0(n29586), .Y(n29588) );
  NAND2XL U33040 ( .A(n29588), .B(n35859), .Y(n15201) );
  AOI32XL U33041 ( .A0(conv_2[11]), .A1(n29590), .A2(n29589), .B0(n33571), 
        .B1(n29590), .Y(n29592) );
  AOI211XL U33042 ( .A0(n29594), .A1(n29592), .B0(n16654), .C0(n29591), .Y(
        n29593) );
  AOI2BB1XL U33043 ( .A0N(n29594), .A1N(n30958), .B0(n29593), .Y(n29595) );
  NAND2XL U33044 ( .A(n29595), .B(n35859), .Y(n15196) );
  OAI2BB1XL U33045 ( .A0N(n29597), .A1N(n29596), .B0(n32876), .Y(n30931) );
  AOI21XL U33046 ( .A0(n29598), .A1(conv_2[235]), .B0(n32876), .Y(n30932) );
  AOI22XL U33047 ( .A0(n33822), .A1(n29600), .B0(conv_2[237]), .B1(n29599), 
        .Y(n29601) );
  NAND2XL U33048 ( .A(n29601), .B(n35859), .Y(n15046) );
  ADDFXL U33049 ( .A(conv_2[216]), .B(n33770), .CI(n29602), .CO(n30155), .S(
        n29603) );
  AOI22XL U33050 ( .A0(n32656), .A1(n29603), .B0(conv_2[216]), .B1(n33765), 
        .Y(n29604) );
  NAND2XL U33051 ( .A(n29604), .B(n35859), .Y(n15062) );
  AOI22XL U33052 ( .A0(n16657), .A1(n29608), .B0(conv_2[206]), .B1(n29607), 
        .Y(n29609) );
  NAND2XL U33053 ( .A(n29609), .B(n35859), .Y(n15067) );
  OAI21XL U33054 ( .A0(n35995), .A1(n29611), .B0(n29610), .Y(n29613) );
  AOI211XL U33055 ( .A0(n29615), .A1(n29613), .B0(n16655), .C0(n29612), .Y(
        n29614) );
  AOI2BB1XL U33056 ( .A0N(n29615), .A1N(n36003), .B0(n29614), .Y(n29616) );
  NAND2XL U33057 ( .A(n29616), .B(n35859), .Y(n14978) );
  NAND2BXL U33058 ( .AN(n29618), .B(n29617), .Y(n29620) );
  AOI211XL U33059 ( .A0(n29622), .A1(n29620), .B0(n16655), .C0(n29619), .Y(
        n29621) );
  AOI2BB1XL U33060 ( .A0N(n29622), .A1N(n35865), .B0(n29621), .Y(n29623) );
  NAND2XL U33061 ( .A(n29623), .B(n35859), .Y(n15177) );
  INVXL U33062 ( .A(conv_2[531]), .Y(n29629) );
  NAND2XL U33063 ( .A(n33629), .B(n29625), .Y(n29624) );
  OAI21XL U33064 ( .A0(n33629), .A1(n29625), .B0(n29624), .Y(n29627) );
  AOI211XL U33065 ( .A0(n29629), .A1(n29627), .B0(n36001), .C0(n29626), .Y(
        n29628) );
  AOI2BB1XL U33066 ( .A0N(n29629), .A1N(n34496), .B0(n29628), .Y(n29630) );
  NAND2XL U33067 ( .A(n29630), .B(n35859), .Y(n14852) );
  INVXL U33068 ( .A(conv_3[498]), .Y(n29636) );
  NAND2XL U33069 ( .A(conv_3[498]), .B(n29634), .Y(n29633) );
  OAI211XL U33070 ( .A0(conv_3[498]), .A1(n29634), .B0(n32660), .C0(n29633), 
        .Y(n29635) );
  OAI211XL U33071 ( .A0(n35841), .A1(n29636), .B0(n35574), .C0(n29635), .Y(
        n15782) );
  NAND2XL U33072 ( .A(conv_3[93]), .B(n29640), .Y(n29639) );
  OAI211XL U33073 ( .A0(conv_3[93]), .A1(n29640), .B0(n31735), .C0(n29639), 
        .Y(n29641) );
  OAI211XL U33074 ( .A0(n35618), .A1(n29642), .B0(n35574), .C0(n29641), .Y(
        n15809) );
  INVXL U33075 ( .A(conv_2[513]), .Y(n29649) );
  AOI21XL U33076 ( .A0(n29645), .A1(n29644), .B0(n29643), .Y(n29647) );
  NAND2XL U33077 ( .A(conv_2[513]), .B(n29647), .Y(n29646) );
  OAI211XL U33078 ( .A0(conv_2[513]), .A1(n29647), .B0(n33778), .C0(n29646), 
        .Y(n29648) );
  OAI211XL U33079 ( .A0(n31013), .A1(n29649), .B0(n34105), .C0(n29648), .Y(
        n15241) );
  NOR2BXL U33080 ( .AN(n29651), .B(n29650), .Y(n29653) );
  NAND2XL U33081 ( .A(conv_3[108]), .B(n29653), .Y(n29652) );
  OAI211XL U33082 ( .A0(conv_3[108]), .A1(n29653), .B0(n24378), .C0(n29652), 
        .Y(n29654) );
  OAI211XL U33083 ( .A0(n34200), .A1(n29655), .B0(n35574), .C0(n29654), .Y(
        n15808) );
  AOI21XL U33084 ( .A0(n29658), .A1(n29657), .B0(n29656), .Y(n29660) );
  NAND2XL U33085 ( .A(conv_3[243]), .B(n29660), .Y(n29659) );
  OAI211XL U33086 ( .A0(conv_3[243]), .A1(n29660), .B0(n30090), .C0(n29659), 
        .Y(n29661) );
  OAI211XL U33087 ( .A0(n35706), .A1(n29662), .B0(n35574), .C0(n29661), .Y(
        n15799) );
  NOR2BXL U33088 ( .AN(n29664), .B(n29663), .Y(n29666) );
  NAND2XL U33089 ( .A(conv_3[34]), .B(n29666), .Y(n29665) );
  OAI211XL U33090 ( .A0(conv_3[34]), .A1(n29666), .B0(n33778), .C0(n29665), 
        .Y(n29667) );
  OAI211XL U33091 ( .A0(n35594), .A1(n29668), .B0(n34097), .C0(n29667), .Y(
        n15777) );
  NAND2XL U33092 ( .A(conv_3[228]), .B(n29672), .Y(n29671) );
  OAI211XL U33093 ( .A0(conv_3[228]), .A1(n29672), .B0(n32052), .C0(n29671), 
        .Y(n29673) );
  OAI211XL U33094 ( .A0(n35676), .A1(n29674), .B0(n35574), .C0(n29673), .Y(
        n15800) );
  NAND2XL U33095 ( .A(n29677), .B(n34768), .Y(n29684) );
  NAND2XL U33096 ( .A(n29678), .B(conv_3[420]), .Y(n29681) );
  INVXL U33097 ( .A(n29681), .Y(n29758) );
  NAND2XL U33098 ( .A(n29679), .B(n29758), .Y(n29682) );
  AOI221XL U33099 ( .A0(n30536), .A1(n29681), .B0(n29680), .B1(n29758), .C0(
        n35499), .Y(n31043) );
  NAND2XL U33100 ( .A(n31043), .B(conv_3[421]), .Y(n31042) );
  NAND2XL U33101 ( .A(n29682), .B(n31042), .Y(n30805) );
  AOI222XL U33102 ( .A0(n30806), .A1(conv_3[422]), .B0(n30806), .B1(n30805), 
        .C0(conv_3[422]), .C1(n30805), .Y(n29683) );
  NAND2XL U33103 ( .A(conv_3[423]), .B(n29686), .Y(n29685) );
  OAI211XL U33104 ( .A0(conv_3[423]), .A1(n29686), .B0(n33712), .C0(n29685), 
        .Y(n29687) );
  OAI211XL U33105 ( .A0(n35778), .A1(n29688), .B0(n35574), .C0(n29687), .Y(
        n15787) );
  INVXL U33106 ( .A(conv_3[198]), .Y(n29694) );
  NOR2BXL U33107 ( .AN(n29690), .B(n29689), .Y(n29692) );
  NAND2XL U33108 ( .A(conv_3[198]), .B(n29692), .Y(n29691) );
  OAI211XL U33109 ( .A0(conv_3[198]), .A1(n29692), .B0(n32656), .C0(n29691), 
        .Y(n29693) );
  OAI211XL U33110 ( .A0(n35646), .A1(n29694), .B0(n35574), .C0(n29693), .Y(
        n15802) );
  INVXL U33111 ( .A(conv_3[393]), .Y(n29700) );
  NAND2XL U33112 ( .A(conv_3[393]), .B(n29698), .Y(n29697) );
  OAI211XL U33113 ( .A0(conv_3[393]), .A1(n29698), .B0(n33712), .C0(n29697), 
        .Y(n29699) );
  OAI211XL U33114 ( .A0(n33703), .A1(n29700), .B0(n35574), .C0(n29699), .Y(
        n15789) );
  INVXL U33115 ( .A(conv_2[34]), .Y(n29706) );
  NAND2XL U33116 ( .A(conv_2[34]), .B(n29704), .Y(n29703) );
  OAI211XL U33117 ( .A0(conv_2[34]), .A1(n29704), .B0(n32660), .C0(n29703), 
        .Y(n29705) );
  OAI211XL U33118 ( .A0(n35865), .A1(n29706), .B0(n34408), .C0(n29705), .Y(
        n15237) );
  INVXL U33119 ( .A(conv_3[438]), .Y(n29712) );
  NOR2BXL U33120 ( .AN(n29708), .B(n29707), .Y(n29710) );
  NAND2XL U33121 ( .A(conv_3[438]), .B(n29710), .Y(n29709) );
  OAI211XL U33122 ( .A0(conv_3[438]), .A1(n29710), .B0(n33712), .C0(n29709), 
        .Y(n29711) );
  OAI211XL U33123 ( .A0(n35792), .A1(n29712), .B0(n35574), .C0(n29711), .Y(
        n15786) );
  NAND2XL U33124 ( .A(conv_2[19]), .B(n29716), .Y(n29715) );
  OAI211XL U33125 ( .A0(conv_2[19]), .A1(n29716), .B0(n32660), .C0(n29715), 
        .Y(n29717) );
  OAI211XL U33126 ( .A0(n30412), .A1(n29718), .B0(n34408), .C0(n29717), .Y(
        n15238) );
  INVXL U33127 ( .A(conv_3[48]), .Y(n29724) );
  XOR2XL U33128 ( .A(n29720), .B(n29719), .Y(n29722) );
  NAND2XL U33129 ( .A(conv_3[48]), .B(n29722), .Y(n29721) );
  OAI211XL U33130 ( .A0(conv_3[48]), .A1(n29722), .B0(n24378), .C0(n29721), 
        .Y(n29723) );
  OAI211XL U33131 ( .A0(n34392), .A1(n29724), .B0(n35574), .C0(n29723), .Y(
        n15812) );
  INVXL U33132 ( .A(conv_3[33]), .Y(n29730) );
  XOR2XL U33133 ( .A(n29726), .B(n29725), .Y(n29728) );
  NAND2XL U33134 ( .A(conv_3[33]), .B(n29728), .Y(n29727) );
  OAI211XL U33135 ( .A0(conv_3[33]), .A1(n29728), .B0(n33778), .C0(n29727), 
        .Y(n29729) );
  OAI211XL U33136 ( .A0(n35594), .A1(n29730), .B0(n35574), .C0(n29729), .Y(
        n15813) );
  INVXL U33137 ( .A(conv_3[183]), .Y(n29737) );
  AOI21XL U33138 ( .A0(n29733), .A1(n29732), .B0(n29731), .Y(n29735) );
  NAND2XL U33139 ( .A(conv_3[183]), .B(n29735), .Y(n29734) );
  OAI211XL U33140 ( .A0(conv_3[183]), .A1(n29735), .B0(n33982), .C0(n29734), 
        .Y(n29736) );
  OAI211XL U33141 ( .A0(n34704), .A1(n29737), .B0(n35574), .C0(n29736), .Y(
        n15803) );
  INVXL U33142 ( .A(conv_2[49]), .Y(n29744) );
  AOI21XL U33143 ( .A0(n29740), .A1(n29739), .B0(n29738), .Y(n29742) );
  NAND2XL U33144 ( .A(conv_2[49]), .B(n29742), .Y(n29741) );
  OAI211XL U33145 ( .A0(conv_2[49]), .A1(n29742), .B0(n32052), .C0(n29741), 
        .Y(n29743) );
  OAI211XL U33146 ( .A0(n34505), .A1(n29744), .B0(n34408), .C0(n29743), .Y(
        n15236) );
  NAND2XL U33147 ( .A(conv_3[156]), .B(n32309), .Y(n32249) );
  NAND2XL U33148 ( .A(n32252), .B(n32249), .Y(n29748) );
  AOI31XL U33149 ( .A0(n36020), .A1(n32248), .A2(n29748), .B0(n16653), .Y(
        n29751) );
  AOI32XL U33150 ( .A0(n32249), .A1(n36020), .A2(n32252), .B0(n29749), .B1(
        n36020), .Y(n29750) );
  INVXL U33151 ( .A(conv_3[157]), .Y(n32250) );
  AOI32XL U33152 ( .A0(n34751), .A1(n29751), .A2(n29750), .B0(n32250), .B1(
        n29751), .Y(n15641) );
  NAND4XL U33153 ( .A(conv_1[56]), .B(conv_1[57]), .C(n35309), .D(n32517), .Y(
        n33050) );
  AND2XL U33154 ( .A(n29753), .B(n29752), .Y(n29754) );
  NOR2X1 U33155 ( .A(n29754), .B(n35309), .Y(n32521) );
  NOR2X1 U33156 ( .A(conv_1[57]), .B(n32521), .Y(n32518) );
  NAND2XL U33157 ( .A(n35316), .B(n32518), .Y(n33049) );
  NAND2XL U33158 ( .A(n33050), .B(n33049), .Y(n29756) );
  NAND2XL U33159 ( .A(conv_1[58]), .B(n29756), .Y(n29755) );
  OAI211XL U33160 ( .A0(conv_1[58]), .A1(n29756), .B0(n33982), .C0(n29755), 
        .Y(n29757) );
  OAI211XL U33161 ( .A0(n35319), .A1(n33048), .B0(n34281), .C0(n29757), .Y(
        n16405) );
  AOI32XL U33162 ( .A0(n29758), .A1(n35778), .A2(n34768), .B0(n16654), .B1(
        n35778), .Y(n29759) );
  AOI32XL U33163 ( .A0(n34742), .A1(n29759), .A2(n34768), .B0(conv_3[420]), 
        .B1(n29759), .Y(n29760) );
  NAND2XL U33164 ( .A(n34755), .B(n29760), .Y(n15895) );
  NAND2XL U33165 ( .A(conv_1[347]), .B(n29765), .Y(n29764) );
  OAI211XL U33166 ( .A0(conv_1[347]), .A1(n29765), .B0(n33778), .C0(n29764), 
        .Y(n29766) );
  OAI211XL U33167 ( .A0(n35447), .A1(n29767), .B0(n29766), .C0(n33542), .Y(
        n16116) );
  NAND2XL U33168 ( .A(conv_2[241]), .B(n29772), .Y(n29771) );
  OAI211XL U33169 ( .A0(conv_2[241]), .A1(n29772), .B0(n33778), .C0(n29771), 
        .Y(n29773) );
  OAI211XL U33170 ( .A0(n35945), .A1(n29774), .B0(n29773), .C0(n35847), .Y(
        n15331) );
  NOR2BXL U33171 ( .AN(n29776), .B(n29775), .Y(n29778) );
  NAND2XL U33172 ( .A(conv_2[526]), .B(n29778), .Y(n29777) );
  OAI211XL U33173 ( .A0(conv_2[526]), .A1(n29778), .B0(n33822), .C0(n29777), 
        .Y(n29779) );
  OAI211XL U33174 ( .A0(n34496), .A1(n29780), .B0(n29779), .C0(n35847), .Y(
        n15312) );
  INVXL U33175 ( .A(conv_2[301]), .Y(n29786) );
  NAND2XL U33176 ( .A(n29782), .B(n29781), .Y(n29784) );
  NAND2XL U33177 ( .A(n29786), .B(n29784), .Y(n29783) );
  OAI211XL U33178 ( .A0(n29786), .A1(n29784), .B0(n32611), .C0(n29783), .Y(
        n29785) );
  OAI211XL U33179 ( .A0(n35976), .A1(n29786), .B0(n29785), .C0(n35847), .Y(
        n15327) );
  NAND2XL U33180 ( .A(n29788), .B(n29787), .Y(n29790) );
  NAND2XL U33181 ( .A(n29792), .B(n29790), .Y(n29789) );
  OAI211XL U33182 ( .A0(n29792), .A1(n29790), .B0(n33778), .C0(n29789), .Y(
        n29791) );
  OAI211XL U33183 ( .A0(n34441), .A1(n29792), .B0(n29791), .C0(n35847), .Y(
        n15317) );
  INVXL U33184 ( .A(conv_2[406]), .Y(n29798) );
  NAND2XL U33185 ( .A(n29794), .B(n29793), .Y(n29796) );
  NAND2XL U33186 ( .A(n29798), .B(n29796), .Y(n29795) );
  OAI211XL U33187 ( .A0(n29798), .A1(n29796), .B0(n33982), .C0(n29795), .Y(
        n29797) );
  OAI211XL U33188 ( .A0(n36047), .A1(n29798), .B0(n29797), .C0(n35847), .Y(
        n15320) );
  NAND2XL U33189 ( .A(n29800), .B(n29799), .Y(n29802) );
  NAND2XL U33190 ( .A(n29804), .B(n29802), .Y(n29801) );
  OAI211XL U33191 ( .A0(n29804), .A1(n29802), .B0(n30090), .C0(n29801), .Y(
        n29803) );
  OAI211XL U33192 ( .A0(n31013), .A1(n29804), .B0(n29803), .C0(n35847), .Y(
        n15313) );
  INVXL U33193 ( .A(conv_2[361]), .Y(n29808) );
  OAI211XL U33194 ( .A0(n29806), .A1(conv_2[361]), .B0(n27932), .C0(n29805), 
        .Y(n29807) );
  OAI211XL U33195 ( .A0(n36017), .A1(n29808), .B0(n29807), .C0(n35847), .Y(
        n15323) );
  INVXL U33196 ( .A(conv_2[331]), .Y(n29814) );
  AND2XL U33197 ( .A(n29810), .B(n29809), .Y(n29812) );
  NAND2XL U33198 ( .A(conv_2[331]), .B(n29812), .Y(n29811) );
  OAI211XL U33199 ( .A0(conv_2[331]), .A1(n29812), .B0(n35336), .C0(n29811), 
        .Y(n29813) );
  OAI211XL U33200 ( .A0(n36003), .A1(n29814), .B0(n29813), .C0(n35847), .Y(
        n15325) );
  NOR2BXL U33201 ( .AN(n29816), .B(n29815), .Y(n29818) );
  NAND2XL U33202 ( .A(conv_2[421]), .B(n29818), .Y(n29817) );
  OAI211XL U33203 ( .A0(conv_2[421]), .A1(n29818), .B0(n33788), .C0(n29817), 
        .Y(n29819) );
  OAI211XL U33204 ( .A0(n36053), .A1(n29820), .B0(n29819), .C0(n35847), .Y(
        n15319) );
  AOI32XL U33205 ( .A0(n29824), .A1(n29823), .A2(n29822), .B0(n29821), .B1(
        n32887), .Y(n29826) );
  AOI211XL U33206 ( .A0(n29828), .A1(n29826), .B0(n16655), .C0(n29825), .Y(
        n29827) );
  NAND2XL U33207 ( .A(n29829), .B(n34281), .Y(n15986) );
  NAND2XL U33208 ( .A(conv_2[170]), .B(n29836), .Y(n29835) );
  OAI211XL U33209 ( .A0(conv_2[170]), .A1(n29836), .B0(n32660), .C0(n29835), 
        .Y(n29837) );
  OAI211XL U33210 ( .A0(n34589), .A1(n29838), .B0(n35859), .C0(n29837), .Y(
        n15093) );
  INVXL U33211 ( .A(conv_2[173]), .Y(n29844) );
  AOI21XL U33212 ( .A0(conv_2[172]), .A1(n29846), .B0(n29831), .Y(n29851) );
  INVXL U33213 ( .A(n29831), .Y(n33974) );
  NAND2XL U33214 ( .A(conv_2[173]), .B(n29842), .Y(n29841) );
  OAI211XL U33215 ( .A0(conv_2[173]), .A1(n29842), .B0(n32611), .C0(n29841), 
        .Y(n29843) );
  OAI211XL U33216 ( .A0(n34589), .A1(n29844), .B0(n35859), .C0(n29843), .Y(
        n15090) );
  INVXL U33217 ( .A(conv_2[172]), .Y(n29850) );
  AOI21XL U33218 ( .A0(n29846), .A1(n29831), .B0(n29845), .Y(n29848) );
  NAND2XL U33219 ( .A(conv_2[172]), .B(n29848), .Y(n29847) );
  OAI211XL U33220 ( .A0(conv_2[172]), .A1(n29848), .B0(n33778), .C0(n29847), 
        .Y(n29849) );
  OAI211XL U33221 ( .A0(n34589), .A1(n29850), .B0(n35859), .C0(n29849), .Y(
        n15091) );
  NOR2X1 U33222 ( .A(n29831), .B(n30894), .Y(n30895) );
  AOI21XL U33223 ( .A0(n30894), .A1(n29831), .B0(n30895), .Y(n29854) );
  NAND2XL U33224 ( .A(conv_2[175]), .B(n29854), .Y(n29853) );
  OAI211XL U33225 ( .A0(conv_2[175]), .A1(n29854), .B0(n34666), .C0(n29853), 
        .Y(n29855) );
  OAI211XL U33226 ( .A0(n34589), .A1(n30897), .B0(n35859), .C0(n29855), .Y(
        n15088) );
  INVXL U33227 ( .A(conv_2[158]), .Y(n29861) );
  AOI2BB1XL U33228 ( .A0N(conv_2[157]), .A1N(n29863), .B0(n34623), .Y(n29856)
         );
  AOI2BB1XL U33229 ( .A0N(n34626), .A1N(n29857), .B0(n29856), .Y(n29859) );
  NAND2XL U33230 ( .A(conv_2[158]), .B(n29859), .Y(n29858) );
  OAI211XL U33231 ( .A0(conv_2[158]), .A1(n29859), .B0(n32181), .C0(n29858), 
        .Y(n29860) );
  OAI211XL U33232 ( .A0(n34631), .A1(n29861), .B0(n35859), .C0(n29860), .Y(
        n15100) );
  AOI21XL U33233 ( .A0(n29863), .A1(n34626), .B0(n29862), .Y(n29865) );
  NAND2XL U33234 ( .A(conv_2[157]), .B(n29865), .Y(n29864) );
  OAI211XL U33235 ( .A0(conv_2[157]), .A1(n29865), .B0(n33822), .C0(n29864), 
        .Y(n29866) );
  OAI211XL U33236 ( .A0(n34631), .A1(n29867), .B0(n35859), .C0(n29866), .Y(
        n15101) );
  INVXL U33237 ( .A(conv_2[256]), .Y(n29871) );
  OAI211XL U33238 ( .A0(conv_2[256]), .A1(n29869), .B0(n28751), .C0(n29868), 
        .Y(n29870) );
  OAI211XL U33239 ( .A0(n34601), .A1(n29871), .B0(n29870), .C0(n35847), .Y(
        n15330) );
  NOR2BXL U33240 ( .AN(n29873), .B(n29872), .Y(n29875) );
  NAND2XL U33241 ( .A(conv_2[317]), .B(n29875), .Y(n29874) );
  OAI211XL U33242 ( .A0(conv_2[317]), .A1(n29875), .B0(n34028), .C0(n29874), 
        .Y(n29876) );
  OAI211XL U33243 ( .A0(n35986), .A1(n29877), .B0(n29876), .C0(n34621), .Y(
        n15290) );
  NAND2XL U33244 ( .A(conv_2[347]), .B(n29882), .Y(n29881) );
  OAI211XL U33245 ( .A0(conv_2[347]), .A1(n29882), .B0(n32660), .C0(n29881), 
        .Y(n29883) );
  OAI211XL U33246 ( .A0(n36010), .A1(n29884), .B0(n29883), .C0(n34621), .Y(
        n15288) );
  AOI21XL U33247 ( .A0(n30946), .A1(n29886), .B0(n29885), .Y(n29888) );
  NAND2XL U33248 ( .A(conv_2[187]), .B(n29888), .Y(n29887) );
  OAI211XL U33249 ( .A0(conv_2[187]), .A1(n29888), .B0(n32656), .C0(n29887), 
        .Y(n29889) );
  OAI211XL U33250 ( .A0(n35917), .A1(n29890), .B0(n35859), .C0(n29889), .Y(
        n15081) );
  NOR2X1 U33251 ( .A(n29891), .B(n30946), .Y(n33455) );
  NOR2X1 U33252 ( .A(conv_2[190]), .B(n33455), .Y(n33456) );
  NOR2X1 U33253 ( .A(n33456), .B(n30946), .Y(n29904) );
  AOI21XL U33254 ( .A0(conv_2[190]), .A1(n33457), .B0(n35914), .Y(n29903) );
  NOR2X1 U33255 ( .A(n30948), .B(n29903), .Y(n30947) );
  NAND3XL U33256 ( .A(n30947), .B(conv_2[192]), .C(n30946), .Y(n29954) );
  INVXL U33257 ( .A(conv_2[192]), .Y(n30952) );
  NAND3XL U33258 ( .A(n30948), .B(n35914), .C(n30952), .Y(n29953) );
  NAND2XL U33259 ( .A(n29954), .B(n29953), .Y(n29895) );
  NAND2XL U33260 ( .A(conv_2[193]), .B(n29895), .Y(n29894) );
  OAI211XL U33261 ( .A0(conv_2[193]), .A1(n29895), .B0(n16657), .C0(n29894), 
        .Y(n29896) );
  OAI211XL U33262 ( .A0(n35917), .A1(n29952), .B0(n35859), .C0(n29896), .Y(
        n15075) );
  NAND2XL U33263 ( .A(conv_2[185]), .B(n29900), .Y(n29899) );
  OAI211XL U33264 ( .A0(conv_2[185]), .A1(n29900), .B0(n16657), .C0(n29899), 
        .Y(n29901) );
  OAI211XL U33265 ( .A0(n35917), .A1(n29902), .B0(n35859), .C0(n29901), .Y(
        n15083) );
  NAND2XL U33266 ( .A(conv_2[191]), .B(n29906), .Y(n29905) );
  OAI211XL U33267 ( .A0(conv_2[191]), .A1(n29906), .B0(n16657), .C0(n29905), 
        .Y(n29907) );
  OAI211XL U33268 ( .A0(n35917), .A1(n29908), .B0(n35859), .C0(n29907), .Y(
        n15077) );
  AOI2BB1XL U33269 ( .A0N(n35914), .A1N(n29910), .B0(n29909), .Y(n29912) );
  NAND2XL U33270 ( .A(conv_2[186]), .B(n29912), .Y(n29911) );
  OAI211XL U33271 ( .A0(conv_2[186]), .A1(n29912), .B0(n16657), .C0(n29911), 
        .Y(n29913) );
  OAI211XL U33272 ( .A0(n35917), .A1(n29914), .B0(n35859), .C0(n29913), .Y(
        n15082) );
  INVXL U33273 ( .A(conv_2[215]), .Y(n29920) );
  NAND2XL U33274 ( .A(conv_2[215]), .B(n29918), .Y(n29917) );
  OAI211XL U33275 ( .A0(conv_2[215]), .A1(n29918), .B0(n33822), .C0(n29917), 
        .Y(n29919) );
  OAI211XL U33276 ( .A0(n35934), .A1(n29920), .B0(n35859), .C0(n29919), .Y(
        n15063) );
  INVXL U33277 ( .A(conv_2[207]), .Y(n29926) );
  AOI21XL U33278 ( .A0(n31310), .A1(n29935), .B0(n29922), .Y(n29924) );
  NAND2XL U33279 ( .A(conv_2[207]), .B(n29924), .Y(n29923) );
  OAI211XL U33280 ( .A0(conv_2[207]), .A1(n29924), .B0(n34028), .C0(n29923), 
        .Y(n29925) );
  OAI211XL U33281 ( .A0(n35931), .A1(n29926), .B0(n35859), .C0(n29925), .Y(
        n15066) );
  AOI2BB1XL U33282 ( .A0N(n29935), .A1N(n29928), .B0(n29927), .Y(n29930) );
  NAND2XL U33283 ( .A(conv_2[204]), .B(n29930), .Y(n29929) );
  OAI211XL U33284 ( .A0(conv_2[204]), .A1(n29930), .B0(n31735), .C0(n29929), 
        .Y(n29931) );
  OAI211XL U33285 ( .A0(n35931), .A1(n29932), .B0(n35859), .C0(n29931), .Y(
        n15069) );
  AOI2BB1XL U33286 ( .A0N(n29935), .A1N(n29934), .B0(n29933), .Y(n29937) );
  NAND2XL U33287 ( .A(conv_2[202]), .B(n29937), .Y(n29936) );
  OAI211XL U33288 ( .A0(conv_2[202]), .A1(n29937), .B0(n16657), .C0(n29936), 
        .Y(n29938) );
  OAI211XL U33289 ( .A0(n35931), .A1(n29939), .B0(n35859), .C0(n29938), .Y(
        n15071) );
  NOR2BXL U33290 ( .AN(n29941), .B(n29940), .Y(n29943) );
  NAND2XL U33291 ( .A(conv_2[200]), .B(n29943), .Y(n29942) );
  OAI211XL U33292 ( .A0(conv_2[200]), .A1(n29943), .B0(n16657), .C0(n29942), 
        .Y(n29944) );
  OAI211XL U33293 ( .A0(n35931), .A1(n29945), .B0(n35859), .C0(n29944), .Y(
        n15073) );
  INVXL U33294 ( .A(conv_2[308]), .Y(n29951) );
  AOI2BB1XL U33295 ( .A0N(n33979), .A1N(n29947), .B0(n29946), .Y(n29949) );
  NAND2XL U33296 ( .A(conv_2[308]), .B(n29949), .Y(n29948) );
  OAI211XL U33297 ( .A0(conv_2[308]), .A1(n29949), .B0(n32052), .C0(n29948), 
        .Y(n29950) );
  OAI211XL U33298 ( .A0(n35976), .A1(n29951), .B0(n34669), .C0(n29950), .Y(
        n15000) );
  AOI22XL U33299 ( .A0(conv_2[193]), .A1(n29954), .B0(n29953), .B1(n29952), 
        .Y(n29956) );
  NAND2XL U33300 ( .A(conv_2[194]), .B(n29956), .Y(n29955) );
  OAI211XL U33301 ( .A0(conv_2[194]), .A1(n29956), .B0(n16657), .C0(n29955), 
        .Y(n29957) );
  OAI211XL U33302 ( .A0(n33442), .A1(n29958), .B0(n35859), .C0(n29957), .Y(
        n15074) );
  INVXL U33303 ( .A(conv_3[153]), .Y(n29964) );
  NOR2BXL U33304 ( .AN(n29960), .B(n29959), .Y(n29962) );
  NAND2XL U33305 ( .A(conv_3[153]), .B(n29962), .Y(n29961) );
  OAI211XL U33306 ( .A0(conv_3[153]), .A1(n29962), .B0(n34028), .C0(n29961), 
        .Y(n29963) );
  OAI211XL U33307 ( .A0(n34751), .A1(n29964), .B0(n35574), .C0(n29963), .Y(
        n15805) );
  INVXL U33308 ( .A(conv_2[407]), .Y(n29970) );
  XOR2XL U33309 ( .A(n29966), .B(n29965), .Y(n29968) );
  NAND2XL U33310 ( .A(conv_2[407]), .B(n29968), .Y(n29967) );
  OAI211XL U33311 ( .A0(conv_2[407]), .A1(n29968), .B0(n33712), .C0(n29967), 
        .Y(n29969) );
  OAI211XL U33312 ( .A0(n36047), .A1(n29970), .B0(n29969), .C0(n34621), .Y(
        n15284) );
  NAND2XL U33313 ( .A(conv_1[486]), .B(n35527), .Y(n35533) );
  NAND2XL U33314 ( .A(conv_1[488]), .B(n35540), .Y(n29983) );
  AOI21XL U33315 ( .A0(conv_1[490]), .A1(n29993), .B0(n35541), .Y(n33209) );
  NAND2XL U33316 ( .A(conv_1[491]), .B(n29975), .Y(n29974) );
  OAI211XL U33317 ( .A0(conv_1[491]), .A1(n29975), .B0(n27932), .C0(n29974), 
        .Y(n29976) );
  OAI211XL U33318 ( .A0(n35544), .A1(n33208), .B0(n16652), .C0(n29976), .Y(
        n15972) );
  ADDFXL U33319 ( .A(conv_3[18]), .B(n29978), .CI(n29977), .CO(n29431), .S(
        n29979) );
  NAND2XL U33320 ( .A(n32656), .B(n29979), .Y(n29980) );
  OAI211XL U33321 ( .A0(n35576), .A1(n29981), .B0(n29980), .C0(n35574), .Y(
        n15814) );
  AOI21XL U33322 ( .A0(n35534), .A1(n29983), .B0(n29982), .Y(n29985) );
  NAND2XL U33323 ( .A(conv_1[489]), .B(n29985), .Y(n29984) );
  OAI211XL U33324 ( .A0(conv_1[489]), .A1(n29985), .B0(n33778), .C0(n29984), 
        .Y(n29986) );
  OAI211XL U33325 ( .A0(n35544), .A1(n29987), .B0(n16652), .C0(n29986), .Y(
        n15974) );
  INVXL U33326 ( .A(conv_2[362]), .Y(n29991) );
  OAI211XL U33327 ( .A0(n29989), .A1(conv_2[362]), .B0(n33982), .C0(n29988), 
        .Y(n29990) );
  OAI211XL U33328 ( .A0(n36017), .A1(n29991), .B0(n29990), .C0(n34621), .Y(
        n15287) );
  INVXL U33329 ( .A(conv_1[490]), .Y(n29997) );
  AOI2BB1XL U33330 ( .A0N(n35541), .A1N(n29993), .B0(n29992), .Y(n29995) );
  NAND2XL U33331 ( .A(conv_1[490]), .B(n29995), .Y(n29994) );
  OAI211XL U33332 ( .A0(conv_1[490]), .A1(n29995), .B0(n34666), .C0(n29994), 
        .Y(n29996) );
  OAI211XL U33333 ( .A0(n35544), .A1(n29997), .B0(n16652), .C0(n29996), .Y(
        n15973) );
  INVXL U33334 ( .A(conv_2[332]), .Y(n30001) );
  NAND2XL U33335 ( .A(conv_2[332]), .B(n29999), .Y(n29998) );
  OAI211XL U33336 ( .A0(conv_2[332]), .A1(n29999), .B0(n33712), .C0(n29998), 
        .Y(n30000) );
  OAI211XL U33337 ( .A0(n36003), .A1(n30001), .B0(n30000), .C0(n34621), .Y(
        n15289) );
  INVXL U33338 ( .A(conv_2[122]), .Y(n30005) );
  NAND2XL U33339 ( .A(conv_2[122]), .B(n30003), .Y(n30002) );
  OAI211XL U33340 ( .A0(conv_2[122]), .A1(n30003), .B0(n16657), .C0(n30002), 
        .Y(n30004) );
  OAI211XL U33341 ( .A0(n34491), .A1(n30005), .B0(n30004), .C0(n34621), .Y(
        n15303) );
  INVXL U33342 ( .A(conv_2[92]), .Y(n30009) );
  NAND2XL U33343 ( .A(conv_2[92]), .B(n30007), .Y(n30006) );
  OAI211XL U33344 ( .A0(conv_2[92]), .A1(n30007), .B0(n34028), .C0(n30006), 
        .Y(n30008) );
  OAI211XL U33345 ( .A0(n34447), .A1(n30009), .B0(n30008), .C0(n34621), .Y(
        n15305) );
  INVXL U33346 ( .A(conv_2[422]), .Y(n30013) );
  NAND2XL U33347 ( .A(conv_2[422]), .B(n30011), .Y(n30010) );
  OAI211XL U33348 ( .A0(conv_2[422]), .A1(n30011), .B0(n33822), .C0(n30010), 
        .Y(n30012) );
  OAI211XL U33349 ( .A0(n36053), .A1(n30013), .B0(n30012), .C0(n34621), .Y(
        n15283) );
  NAND2XL U33350 ( .A(conv_2[452]), .B(n30015), .Y(n30014) );
  OAI211XL U33351 ( .A0(conv_2[452]), .A1(n30015), .B0(n28751), .C0(n30014), 
        .Y(n30016) );
  OAI211XL U33352 ( .A0(n34441), .A1(n30017), .B0(n30016), .C0(n34621), .Y(
        n15281) );
  AOI2BB1XL U33353 ( .A0N(n30044), .A1N(n30019), .B0(n30018), .Y(n30021) );
  NAND2XL U33354 ( .A(conv_1[456]), .B(n30021), .Y(n30020) );
  OAI211XL U33355 ( .A0(conv_1[456]), .A1(n30021), .B0(n33778), .C0(n30020), 
        .Y(n30022) );
  OAI211XL U33356 ( .A0(n30056), .A1(n30023), .B0(n34281), .C0(n30022), .Y(
        n16007) );
  OAI2BB1XL U33357 ( .A0N(n30044), .A1N(n30025), .B0(n30024), .Y(n30027) );
  NAND2XL U33358 ( .A(n30029), .B(n30027), .Y(n30026) );
  OAI211XL U33359 ( .A0(n30029), .A1(n30027), .B0(n33778), .C0(n30026), .Y(
        n30028) );
  OAI211XL U33360 ( .A0(n30056), .A1(n30029), .B0(n16652), .C0(n30028), .Y(
        n16002) );
  NAND2XL U33361 ( .A(conv_1[459]), .B(n30033), .Y(n30032) );
  OAI211XL U33362 ( .A0(conv_1[459]), .A1(n30033), .B0(n32660), .C0(n30032), 
        .Y(n30034) );
  OAI211XL U33363 ( .A0(n30056), .A1(n30035), .B0(n34689), .C0(n30034), .Y(
        n16004) );
  AOI2BB1XL U33364 ( .A0N(n30044), .A1N(n30037), .B0(n30036), .Y(n30039) );
  NAND2XL U33365 ( .A(conv_1[458]), .B(n30039), .Y(n30038) );
  OAI211XL U33366 ( .A0(conv_1[458]), .A1(n30039), .B0(n33778), .C0(n30038), 
        .Y(n30040) );
  OAI211XL U33367 ( .A0(n30056), .A1(n30041), .B0(n34544), .C0(n30040), .Y(
        n16005) );
  OAI21XL U33368 ( .A0(n30044), .A1(n30043), .B0(n30042), .Y(n30046) );
  NAND2XL U33369 ( .A(n30048), .B(n30046), .Y(n30045) );
  OAI211XL U33370 ( .A0(n30048), .A1(n30046), .B0(n33982), .C0(n30045), .Y(
        n30047) );
  OAI211XL U33371 ( .A0(n30056), .A1(n30048), .B0(n34544), .C0(n30047), .Y(
        n16003) );
  AOI21XL U33372 ( .A0(n30051), .A1(n30050), .B0(n30049), .Y(n30053) );
  NAND2XL U33373 ( .A(conv_1[457]), .B(n30053), .Y(n30052) );
  OAI211XL U33374 ( .A0(conv_1[457]), .A1(n30053), .B0(n33778), .C0(n30052), 
        .Y(n30054) );
  OAI211XL U33375 ( .A0(n30056), .A1(n30055), .B0(n34682), .C0(n30054), .Y(
        n16006) );
  INVXL U33376 ( .A(conv_1[360]), .Y(n30060) );
  OAI211XL U33377 ( .A0(conv_1[360]), .A1(n30058), .B0(n33778), .C0(n30057), 
        .Y(n30059) );
  OAI211XL U33378 ( .A0(n35458), .A1(n30060), .B0(n30059), .C0(n34773), .Y(
        n16103) );
  NAND2XL U33379 ( .A(conv_2[127]), .B(n30064), .Y(n30063) );
  OAI211XL U33380 ( .A0(conv_2[127]), .A1(n30064), .B0(n16657), .C0(n30063), 
        .Y(n30065) );
  OAI211XL U33381 ( .A0(n34491), .A1(n30066), .B0(n33815), .C0(n30065), .Y(
        n15121) );
  INVXL U33382 ( .A(conv_2[133]), .Y(n30441) );
  NAND2XL U33383 ( .A(n30444), .B(n30443), .Y(n30442) );
  OAI21XL U33384 ( .A0(n30444), .A1(n30443), .B0(n30442), .Y(n30069) );
  NAND2XL U33385 ( .A(conv_2[133]), .B(n30069), .Y(n30068) );
  OAI211XL U33386 ( .A0(conv_2[133]), .A1(n30069), .B0(n30090), .C0(n30068), 
        .Y(n30070) );
  OAI211XL U33387 ( .A0(n34491), .A1(n30441), .B0(n33815), .C0(n30070), .Y(
        n15115) );
  OAI32XL U33388 ( .A0(n30443), .A1(conv_2[129]), .A2(n34343), .B0(n34344), 
        .B1(n30071), .Y(n30073) );
  NAND2XL U33389 ( .A(conv_2[130]), .B(n30073), .Y(n30072) );
  OAI211XL U33390 ( .A0(conv_2[130]), .A1(n30073), .B0(n30090), .C0(n30072), 
        .Y(n30074) );
  OAI211XL U33391 ( .A0(n34491), .A1(n30075), .B0(n33815), .C0(n30074), .Y(
        n15118) );
  INVXL U33392 ( .A(conv_2[141]), .Y(n30081) );
  AOI2BB1XL U33393 ( .A0N(n35907), .A1N(n30077), .B0(n30076), .Y(n30079) );
  NAND2XL U33394 ( .A(conv_2[141]), .B(n30079), .Y(n30078) );
  OAI211XL U33395 ( .A0(conv_2[141]), .A1(n30079), .B0(n30090), .C0(n30078), 
        .Y(n30080) );
  OAI211XL U33396 ( .A0(n35902), .A1(n30081), .B0(n33815), .C0(n30080), .Y(
        n15112) );
  AOI32XL U33397 ( .A0(conv_2[146]), .A1(n30082), .A2(n34357), .B0(n35907), 
        .B1(n30082), .Y(n30084) );
  NAND2XL U33398 ( .A(n30086), .B(n30084), .Y(n30083) );
  OAI211XL U33399 ( .A0(n30086), .A1(n30084), .B0(n33778), .C0(n30083), .Y(
        n30085) );
  OAI211XL U33400 ( .A0(n35902), .A1(n30086), .B0(n33815), .C0(n30085), .Y(
        n15106) );
  AOI21XL U33401 ( .A0(n35899), .A1(n30088), .B0(n30087), .Y(n30091) );
  NAND2XL U33402 ( .A(conv_2[144]), .B(n30091), .Y(n30089) );
  OAI211XL U33403 ( .A0(conv_2[144]), .A1(n30091), .B0(n30090), .C0(n30089), 
        .Y(n30092) );
  OAI211XL U33404 ( .A0(n35902), .A1(n30093), .B0(n33815), .C0(n30092), .Y(
        n15109) );
  AOI2BB1XL U33405 ( .A0N(n35907), .A1N(n30095), .B0(n30094), .Y(n30097) );
  NAND2XL U33406 ( .A(conv_2[145]), .B(n30097), .Y(n30096) );
  OAI211XL U33407 ( .A0(conv_2[145]), .A1(n30097), .B0(n32611), .C0(n30096), 
        .Y(n30098) );
  OAI211XL U33408 ( .A0(n35902), .A1(n30099), .B0(n33815), .C0(n30098), .Y(
        n15108) );
  AOI21XL U33409 ( .A0(n30242), .A1(n30101), .B0(n30100), .Y(n30103) );
  NAND2XL U33410 ( .A(conv_2[66]), .B(n30103), .Y(n30102) );
  OAI211XL U33411 ( .A0(conv_2[66]), .A1(n30103), .B0(n16657), .C0(n30102), 
        .Y(n30104) );
  OAI211XL U33412 ( .A0(n35846), .A1(n30105), .B0(n33815), .C0(n30104), .Y(
        n15162) );
  AOI21XL U33413 ( .A0(conv_2[67]), .A1(n30107), .B0(n33735), .Y(n30119) );
  NAND2XL U33414 ( .A(conv_2[68]), .B(n30109), .Y(n30108) );
  OAI211XL U33415 ( .A0(conv_2[68]), .A1(n30109), .B0(n16657), .C0(n30108), 
        .Y(n30110) );
  OAI211XL U33416 ( .A0(n35846), .A1(n30111), .B0(n33815), .C0(n30110), .Y(
        n15160) );
  INVXL U33417 ( .A(conv_2[65]), .Y(n30117) );
  NOR2BXL U33418 ( .AN(n30113), .B(n30112), .Y(n30115) );
  NAND2XL U33419 ( .A(conv_2[65]), .B(n30115), .Y(n30114) );
  OAI211XL U33420 ( .A0(conv_2[65]), .A1(n30115), .B0(n16657), .C0(n30114), 
        .Y(n30116) );
  OAI211XL U33421 ( .A0(n35846), .A1(n30117), .B0(n33815), .C0(n30116), .Y(
        n15163) );
  NAND2XL U33422 ( .A(n30977), .B(n30972), .Y(n30125) );
  OAI2BB1XL U33423 ( .A0N(conv_2[69]), .A1N(n30973), .B0(n30242), .Y(n30126)
         );
  OAI2BB1XL U33424 ( .A0N(n33735), .A1N(n30125), .B0(n30126), .Y(n30122) );
  NAND2XL U33425 ( .A(n30124), .B(n30122), .Y(n30121) );
  OAI211XL U33426 ( .A0(n30124), .A1(n30122), .B0(n33788), .C0(n30121), .Y(
        n30123) );
  OAI211XL U33427 ( .A0(n35846), .A1(n30124), .B0(n33815), .C0(n30123), .Y(
        n15158) );
  INVXL U33428 ( .A(conv_2[71]), .Y(n30130) );
  NAND2XL U33429 ( .A(conv_2[71]), .B(n30128), .Y(n30127) );
  OAI211XL U33430 ( .A0(conv_2[71]), .A1(n30128), .B0(n16657), .C0(n30127), 
        .Y(n30129) );
  OAI211XL U33431 ( .A0(n35846), .A1(n30130), .B0(n33815), .C0(n30129), .Y(
        n15157) );
  INVXL U33432 ( .A(conv_1[361]), .Y(n30134) );
  NAND2XL U33433 ( .A(conv_1[361]), .B(n30132), .Y(n30131) );
  OAI211XL U33434 ( .A0(conv_1[361]), .A1(n30132), .B0(n16656), .C0(n30131), 
        .Y(n30133) );
  OAI211XL U33435 ( .A0(n35458), .A1(n30134), .B0(n30133), .C0(n33067), .Y(
        n16102) );
  NAND4XL U33436 ( .A(conv_2[116]), .B(conv_2[117]), .C(n35884), .D(n34642), 
        .Y(n30250) );
  INVXL U33437 ( .A(n35884), .Y(n35891) );
  OAI21XL U33438 ( .A0(conv_2[115]), .A1(n30148), .B0(n35891), .Y(n34643) );
  NAND2XL U33439 ( .A(n34647), .B(n34643), .Y(n30138) );
  NAND3XL U33440 ( .A(n35891), .B(n34368), .C(n34364), .Y(n30249) );
  NAND2XL U33441 ( .A(n30250), .B(n30249), .Y(n30140) );
  NAND2XL U33442 ( .A(conv_2[118]), .B(n30140), .Y(n30139) );
  OAI211XL U33443 ( .A0(conv_2[118]), .A1(n30140), .B0(n33778), .C0(n30139), 
        .Y(n30141) );
  OAI211XL U33444 ( .A0(n35894), .A1(n30248), .B0(n33815), .C0(n30141), .Y(
        n15125) );
  INVXL U33445 ( .A(conv_2[111]), .Y(n30147) );
  OAI2BB1XL U33446 ( .A0N(n35891), .A1N(n30143), .B0(n30142), .Y(n30145) );
  NAND2XL U33447 ( .A(n30147), .B(n30145), .Y(n30144) );
  OAI211XL U33448 ( .A0(n30147), .A1(n30145), .B0(n34028), .C0(n30144), .Y(
        n30146) );
  OAI211XL U33449 ( .A0(n35894), .A1(n30147), .B0(n33815), .C0(n30146), .Y(
        n15132) );
  INVXL U33450 ( .A(conv_2[115]), .Y(n30153) );
  AOI2BB1XL U33451 ( .A0N(n35891), .A1N(n30149), .B0(n30148), .Y(n30151) );
  NAND2XL U33452 ( .A(conv_2[115]), .B(n30151), .Y(n30150) );
  OAI211XL U33453 ( .A0(conv_2[115]), .A1(n30151), .B0(n32181), .C0(n30150), 
        .Y(n30152) );
  OAI211XL U33454 ( .A0(n35894), .A1(n30153), .B0(n33815), .C0(n30152), .Y(
        n15128) );
  AOI21XL U33455 ( .A0(n30155), .A1(n33770), .B0(n30154), .Y(n30157) );
  NAND2XL U33456 ( .A(conv_2[217]), .B(n30157), .Y(n30156) );
  OAI211XL U33457 ( .A0(conv_2[217]), .A1(n30157), .B0(n16657), .C0(n30156), 
        .Y(n30158) );
  OAI211XL U33458 ( .A0(n35934), .A1(n30159), .B0(n33815), .C0(n30158), .Y(
        n15061) );
  INVXL U33459 ( .A(conv_2[57]), .Y(n31136) );
  NAND2XL U33460 ( .A(n30161), .B(n30160), .Y(n30162) );
  AOI32XL U33461 ( .A0(conv_2[56]), .A1(n31135), .A2(n31133), .B0(n31137), 
        .B1(n31135), .Y(n30164) );
  NAND2XL U33462 ( .A(n31136), .B(n30164), .Y(n30163) );
  OAI211XL U33463 ( .A0(n31136), .A1(n30164), .B0(n16657), .C0(n30163), .Y(
        n30165) );
  OAI211XL U33464 ( .A0(n34505), .A1(n31136), .B0(n33815), .C0(n30165), .Y(
        n15166) );
  AOI21XL U33465 ( .A0(n30924), .A1(n30167), .B0(n30166), .Y(n30169) );
  NAND2XL U33466 ( .A(conv_2[82]), .B(n30169), .Y(n30168) );
  OAI211XL U33467 ( .A0(conv_2[82]), .A1(n30169), .B0(n34666), .C0(n30168), 
        .Y(n30170) );
  OAI211XL U33468 ( .A0(n35879), .A1(n30171), .B0(n33815), .C0(n30170), .Y(
        n15151) );
  AOI21XL U33469 ( .A0(conv_2[85]), .A1(n33813), .B0(n35876), .Y(n31002) );
  AOI22XL U33470 ( .A0(n35876), .A1(n30927), .B0(n30925), .B1(n30924), .Y(
        n30176) );
  NAND2XL U33471 ( .A(n30926), .B(n30176), .Y(n30175) );
  OAI211XL U33472 ( .A0(n30926), .A1(n30176), .B0(n34666), .C0(n30175), .Y(
        n30177) );
  OAI211XL U33473 ( .A0(n35879), .A1(n30926), .B0(n33815), .C0(n30177), .Y(
        n15146) );
  NAND2XL U33474 ( .A(conv_2[80]), .B(n30181), .Y(n30180) );
  OAI211XL U33475 ( .A0(conv_2[80]), .A1(n30181), .B0(n34666), .C0(n30180), 
        .Y(n30182) );
  OAI211XL U33476 ( .A0(n35879), .A1(n30183), .B0(n33815), .C0(n30182), .Y(
        n15153) );
  NAND2XL U33477 ( .A(conv_3[468]), .B(n30187), .Y(n30186) );
  OAI211XL U33478 ( .A0(conv_3[468]), .A1(n30187), .B0(n16656), .C0(n30186), 
        .Y(n30188) );
  OAI211XL U33479 ( .A0(n35813), .A1(n30189), .B0(n35574), .C0(n30188), .Y(
        n15784) );
  NAND2XL U33480 ( .A(n32611), .B(n30192), .Y(n30193) );
  OAI211XL U33481 ( .A0(n34080), .A1(n30194), .B0(n34682), .C0(n30193), .Y(
        n16198) );
  OAI31XL U33482 ( .A0(conv_3[21]), .A1(conv_3[22]), .A2(n31274), .B0(n33002), 
        .Y(n31267) );
  INVXL U33483 ( .A(n33002), .Y(n31304) );
  AOI21XL U33484 ( .A0(n31272), .A1(n31267), .B0(n31304), .Y(n30199) );
  INVXL U33485 ( .A(conv_3[22]), .Y(n31266) );
  NAND2XL U33486 ( .A(conv_3[23]), .B(n31268), .Y(n31250) );
  NAND2XL U33487 ( .A(n31304), .B(n31250), .Y(n30198) );
  AOI31XL U33488 ( .A0(n36020), .A1(n31252), .A2(n30198), .B0(n16653), .Y(
        n30201) );
  AOI32XL U33489 ( .A0(n31250), .A1(n36020), .A2(n31304), .B0(n30199), .B1(
        n36020), .Y(n30200) );
  INVXL U33490 ( .A(conv_3[24]), .Y(n31251) );
  AOI32XL U33491 ( .A0(n35576), .A1(n30201), .A2(n30200), .B0(n31251), .B1(
        n30201), .Y(n15729) );
  INVXL U33492 ( .A(conv_2[100]), .Y(n30214) );
  OAI2BB1XL U33493 ( .A0N(n30202), .A1N(conv_2[97]), .B0(n30225), .Y(n30220)
         );
  NAND2XL U33494 ( .A(n30940), .B(n30203), .Y(n30219) );
  NAND2XL U33495 ( .A(n30224), .B(n30219), .Y(n30939) );
  NAND2XL U33496 ( .A(n30214), .B(n30205), .Y(n30206) );
  OAI21XL U33497 ( .A0(conv_2[101]), .A1(n30206), .B0(n30940), .Y(n30227) );
  OAI21XL U33498 ( .A0(n30940), .A1(n30226), .B0(n30227), .Y(n30208) );
  NAND2XL U33499 ( .A(n30228), .B(n30208), .Y(n30207) );
  OAI211XL U33500 ( .A0(n30228), .A1(n30208), .B0(n16657), .C0(n30207), .Y(
        n30209) );
  OAI211XL U33501 ( .A0(n34447), .A1(n30228), .B0(n33815), .C0(n30209), .Y(
        n15136) );
  OAI2BB1XL U33502 ( .A0N(n30212), .A1N(n30214), .B0(n30211), .Y(n30213) );
  OAI211XL U33503 ( .A0(n34447), .A1(n30214), .B0(n33815), .C0(n30213), .Y(
        n15138) );
  OAI2BB1XL U33504 ( .A0N(n30216), .A1N(n30218), .B0(n30215), .Y(n30217) );
  OAI211XL U33505 ( .A0(n34447), .A1(n30218), .B0(n33815), .C0(n30217), .Y(
        n15137) );
  NAND2XL U33506 ( .A(n30220), .B(n30219), .Y(n30222) );
  NAND2XL U33507 ( .A(n30224), .B(n30222), .Y(n30221) );
  OAI211XL U33508 ( .A0(n30224), .A1(n30222), .B0(n33982), .C0(n30221), .Y(
        n30223) );
  OAI211XL U33509 ( .A0(n34447), .A1(n30224), .B0(n33815), .C0(n30223), .Y(
        n15140) );
  NAND3XL U33510 ( .A(n30226), .B(conv_2[102]), .C(n30225), .Y(n33289) );
  NAND3XL U33511 ( .A(n30940), .B(n30228), .C(n30227), .Y(n33288) );
  AOI22XL U33512 ( .A0(conv_2[103]), .A1(n33289), .B0(n33288), .B1(n33292), 
        .Y(n30230) );
  NAND2XL U33513 ( .A(conv_2[104]), .B(n30230), .Y(n30229) );
  OAI211XL U33514 ( .A0(conv_2[104]), .A1(n30230), .B0(n33822), .C0(n30229), 
        .Y(n30231) );
  OAI211XL U33515 ( .A0(n34520), .A1(n30232), .B0(n33815), .C0(n30231), .Y(
        n15134) );
  AOI22XL U33516 ( .A0(conv_2[148]), .A1(n30235), .B0(n30234), .B1(n30233), 
        .Y(n30237) );
  NAND2XL U33517 ( .A(conv_2[149]), .B(n30237), .Y(n30236) );
  OAI211XL U33518 ( .A0(conv_2[149]), .A1(n30237), .B0(n16657), .C0(n30236), 
        .Y(n30238) );
  OAI211XL U33519 ( .A0(n33853), .A1(n30239), .B0(n33815), .C0(n30238), .Y(
        n15104) );
  NOR2X1 U33520 ( .A(conv_2[71]), .B(n30240), .Y(n30243) );
  NAND3XL U33521 ( .A(n33734), .B(conv_2[72]), .C(n30242), .Y(n34725) );
  NAND2XL U33522 ( .A(n33735), .B(n33733), .Y(n34724) );
  INVXL U33523 ( .A(conv_2[73]), .Y(n34728) );
  AOI22XL U33524 ( .A0(conv_2[73]), .A1(n34725), .B0(n34724), .B1(n34728), .Y(
        n30245) );
  NAND2XL U33525 ( .A(conv_2[74]), .B(n30245), .Y(n30244) );
  OAI211XL U33526 ( .A0(conv_2[74]), .A1(n30245), .B0(n34666), .C0(n30244), 
        .Y(n30246) );
  OAI211XL U33527 ( .A0(n34676), .A1(n30247), .B0(n33815), .C0(n30246), .Y(
        n15154) );
  AOI22XL U33528 ( .A0(conv_2[118]), .A1(n30250), .B0(n30249), .B1(n30248), 
        .Y(n30252) );
  NAND2XL U33529 ( .A(conv_2[119]), .B(n30252), .Y(n30251) );
  OAI211XL U33530 ( .A0(conv_2[119]), .A1(n30252), .B0(n33982), .C0(n30251), 
        .Y(n30253) );
  OAI211XL U33531 ( .A0(n34520), .A1(n30254), .B0(n33815), .C0(n30253), .Y(
        n15124) );
  AOI22XL U33532 ( .A0(n32611), .A1(intadd_1_SUM_1_), .B0(conv_1[424]), .B1(
        n35510), .Y(n30255) );
  NAND2XL U33533 ( .A(n30255), .B(n35489), .Y(n16039) );
  NAND2XL U33534 ( .A(n30257), .B(n30256), .Y(n30259) );
  NAND2XL U33535 ( .A(conv_1[523]), .B(n30259), .Y(n30258) );
  OAI211XL U33536 ( .A0(conv_1[523]), .A1(n30259), .B0(n33778), .C0(n30258), 
        .Y(n30260) );
  OAI211XL U33537 ( .A0(n35547), .A1(n30261), .B0(n34281), .C0(n30260), .Y(
        n15940) );
  OAI211XL U33538 ( .A0(n30262), .A1(conv_1[519]), .B0(n34028), .C0(n30266), 
        .Y(n30263) );
  OAI211XL U33539 ( .A0(n35547), .A1(n30264), .B0(n34696), .C0(n30263), .Y(
        n15944) );
  AOI21XL U33540 ( .A0(n30267), .A1(n30266), .B0(n30265), .Y(n30269) );
  NAND2XL U33541 ( .A(conv_1[520]), .B(n30269), .Y(n30268) );
  OAI211XL U33542 ( .A0(conv_1[520]), .A1(n30269), .B0(n33778), .C0(n30268), 
        .Y(n30270) );
  OAI211XL U33543 ( .A0(n35547), .A1(n30271), .B0(n16652), .C0(n30270), .Y(
        n15943) );
  ADDFXL U33544 ( .A(conv_2[242]), .B(n30273), .CI(n30272), .CO(n28145), .S(
        n30274) );
  AOI22XL U33545 ( .A0(n33778), .A1(n30274), .B0(conv_2[242]), .B1(n33679), 
        .Y(n30275) );
  NAND2XL U33546 ( .A(n30275), .B(n34621), .Y(n15295) );
  INVXL U33547 ( .A(conv_1[364]), .Y(n30281) );
  NAND2XL U33548 ( .A(conv_1[364]), .B(n30279), .Y(n30278) );
  OAI211XL U33549 ( .A0(conv_1[364]), .A1(n30279), .B0(n32052), .C0(n30278), 
        .Y(n30280) );
  OAI211XL U33550 ( .A0(n35458), .A1(n30281), .B0(n35489), .C0(n30280), .Y(
        n16099) );
  INVXL U33551 ( .A(conv_1[349]), .Y(n30287) );
  NAND2XL U33552 ( .A(conv_1[349]), .B(n30285), .Y(n30284) );
  OAI211XL U33553 ( .A0(conv_1[349]), .A1(n30285), .B0(n33982), .C0(n30284), 
        .Y(n30286) );
  OAI211XL U33554 ( .A0(n35447), .A1(n30287), .B0(n35489), .C0(n30286), .Y(
        n16114) );
  NAND2XL U33555 ( .A(n30289), .B(n30288), .Y(n30291) );
  NAND2XL U33556 ( .A(n30293), .B(n30291), .Y(n30290) );
  OAI211XL U33557 ( .A0(n30293), .A1(n30291), .B0(n33778), .C0(n30290), .Y(
        n30292) );
  OAI211XL U33558 ( .A0(n34137), .A1(n30293), .B0(n35847), .C0(n30292), .Y(
        n15315) );
  OAI211XL U33559 ( .A0(n30295), .A1(conv_2[466]), .B0(n27932), .C0(n30294), 
        .Y(n30296) );
  OAI211XL U33560 ( .A0(n34177), .A1(n30297), .B0(n35847), .C0(n30296), .Y(
        n15316) );
  INVXL U33561 ( .A(conv_2[376]), .Y(n30301) );
  OAI211XL U33562 ( .A0(n30299), .A1(conv_2[376]), .B0(n33778), .C0(n30298), 
        .Y(n30300) );
  OAI211XL U33563 ( .A0(n36028), .A1(n30301), .B0(n35847), .C0(n30300), .Y(
        n15322) );
  OAI211XL U33564 ( .A0(n30303), .A1(conv_2[286]), .B0(n33778), .C0(n30302), 
        .Y(n30304) );
  OAI211XL U33565 ( .A0(n35963), .A1(n30305), .B0(n35847), .C0(n30304), .Y(
        n15328) );
  INVXL U33566 ( .A(conv_2[391]), .Y(n30311) );
  NOR2BXL U33567 ( .AN(n30307), .B(n30306), .Y(n30309) );
  NAND2XL U33568 ( .A(conv_2[391]), .B(n30309), .Y(n30308) );
  OAI211XL U33569 ( .A0(conv_2[391]), .A1(n30309), .B0(n30090), .C0(n30308), 
        .Y(n30310) );
  OAI211XL U33570 ( .A0(n36031), .A1(n30311), .B0(n35847), .C0(n30310), .Y(
        n15321) );
  INVXL U33571 ( .A(conv_2[436]), .Y(n30317) );
  NOR2BXL U33572 ( .AN(n30313), .B(n30312), .Y(n30315) );
  NAND2XL U33573 ( .A(conv_2[436]), .B(n30315), .Y(n30314) );
  OAI211XL U33574 ( .A0(conv_2[436]), .A1(n30315), .B0(n31735), .C0(n30314), 
        .Y(n30316) );
  OAI211XL U33575 ( .A0(n36070), .A1(n30317), .B0(n35847), .C0(n30316), .Y(
        n15318) );
  NAND2XL U33576 ( .A(conv_2[497]), .B(n30321), .Y(n30320) );
  OAI211XL U33577 ( .A0(conv_2[497]), .A1(n30321), .B0(n33712), .C0(n30320), 
        .Y(n30322) );
  OAI211XL U33578 ( .A0(n36091), .A1(n30323), .B0(n34621), .C0(n30322), .Y(
        n15278) );
  OAI21XL U33579 ( .A0(n33208), .A1(n33209), .B0(n35534), .Y(n30327) );
  AOI31XL U33580 ( .A0(n36020), .A1(n33210), .A2(n30327), .B0(n35549), .Y(
        n30330) );
  INVXL U33581 ( .A(n30326), .Y(n30328) );
  OAI2BB1XL U33582 ( .A0N(n30328), .A1N(n30327), .B0(n35336), .Y(n30329) );
  INVXL U33583 ( .A(conv_1[492]), .Y(n33207) );
  AOI32XL U33584 ( .A0(n35544), .A1(n30330), .A2(n30329), .B0(n33207), .B1(
        n30330), .Y(n15971) );
  XOR2XL U33585 ( .A(n30332), .B(n30331), .Y(n30334) );
  NAND2XL U33586 ( .A(conv_2[467]), .B(n30334), .Y(n30333) );
  OAI211XL U33587 ( .A0(conv_2[467]), .A1(n30334), .B0(n36020), .C0(n30333), 
        .Y(n30335) );
  OAI211XL U33588 ( .A0(n34177), .A1(n30336), .B0(n34621), .C0(n30335), .Y(
        n15280) );
  XOR2XL U33589 ( .A(n30338), .B(n30337), .Y(n30340) );
  NAND2XL U33590 ( .A(conv_2[482]), .B(n30340), .Y(n30339) );
  OAI211XL U33591 ( .A0(conv_2[482]), .A1(n30340), .B0(n34666), .C0(n30339), 
        .Y(n30341) );
  OAI211XL U33592 ( .A0(n34137), .A1(n30342), .B0(n34621), .C0(n30341), .Y(
        n15279) );
  INVXL U33593 ( .A(conv_2[392]), .Y(n30348) );
  NAND2XL U33594 ( .A(conv_2[392]), .B(n30346), .Y(n30345) );
  OAI211XL U33595 ( .A0(conv_2[392]), .A1(n30346), .B0(n33822), .C0(n30345), 
        .Y(n30347) );
  OAI211XL U33596 ( .A0(n36031), .A1(n30348), .B0(n34621), .C0(n30347), .Y(
        n15285) );
  INVXL U33597 ( .A(filter_3[12]), .Y(n30351) );
  INVXL U33598 ( .A(filter_3[6]), .Y(n36101) );
  AOI22XL U33599 ( .A0(n36107), .A1(n30351), .B0(n36101), .B1(n30392), .Y(
        n14742) );
  INVXL U33600 ( .A(filter_3[13]), .Y(n30364) );
  INVXL U33601 ( .A(filter_3[7]), .Y(n36106) );
  AOI22XL U33602 ( .A0(n36107), .A1(n30364), .B0(n36106), .B1(n30392), .Y(
        n14743) );
  INVXL U33603 ( .A(filter_3[14]), .Y(n30352) );
  INVXL U33604 ( .A(filter_3[8]), .Y(n36105) );
  AOI22XL U33605 ( .A0(n36107), .A1(n30352), .B0(n36105), .B1(n30392), .Y(
        n14744) );
  INVXL U33606 ( .A(filter_3[15]), .Y(n30353) );
  INVXL U33607 ( .A(filter_3[9]), .Y(n36104) );
  AOI22XL U33608 ( .A0(n36107), .A1(n30353), .B0(n36104), .B1(n30392), .Y(
        n14745) );
  INVXL U33609 ( .A(filter_3[16]), .Y(n30354) );
  INVXL U33610 ( .A(filter_3[10]), .Y(n36103) );
  AOI22XL U33611 ( .A0(n36107), .A1(n30354), .B0(n36103), .B1(n30392), .Y(
        n14746) );
  INVXL U33612 ( .A(filter_3[17]), .Y(n30355) );
  INVXL U33613 ( .A(filter_3[11]), .Y(n36102) );
  AOI22XL U33614 ( .A0(n36107), .A1(n30355), .B0(n36102), .B1(n30392), .Y(
        n14747) );
  INVXL U33615 ( .A(filter_3[18]), .Y(n30356) );
  AOI22XL U33616 ( .A0(n36107), .A1(n30356), .B0(n30351), .B1(n30392), .Y(
        n14748) );
  INVXL U33617 ( .A(filter_3[20]), .Y(n30357) );
  AOI22XL U33618 ( .A0(n36107), .A1(n30357), .B0(n30352), .B1(n30392), .Y(
        n14750) );
  INVXL U33619 ( .A(filter_3[21]), .Y(n30358) );
  AOI22XL U33620 ( .A0(n36107), .A1(n30358), .B0(n30353), .B1(n30392), .Y(
        n14751) );
  INVXL U33621 ( .A(filter_3[22]), .Y(n30359) );
  AOI22XL U33622 ( .A0(n36107), .A1(n30359), .B0(n30354), .B1(n30392), .Y(
        n14752) );
  INVXL U33623 ( .A(filter_3[23]), .Y(n30360) );
  AOI22XL U33624 ( .A0(n36107), .A1(n30360), .B0(n30355), .B1(n30392), .Y(
        n14753) );
  INVXL U33625 ( .A(filter_3[24]), .Y(n30361) );
  AOI22XL U33626 ( .A0(n36107), .A1(n30361), .B0(n30356), .B1(n30392), .Y(
        n14754) );
  INVXL U33627 ( .A(filter_3[25]), .Y(n30362) );
  INVXL U33628 ( .A(filter_3[19]), .Y(n30365) );
  AOI22XL U33629 ( .A0(n36107), .A1(n30362), .B0(n30365), .B1(n30392), .Y(
        n14755) );
  INVXL U33630 ( .A(filter_3[26]), .Y(n30363) );
  AOI22XL U33631 ( .A0(n36107), .A1(n30363), .B0(n30357), .B1(n30392), .Y(
        n14756) );
  INVXL U33632 ( .A(filter_3[27]), .Y(n30366) );
  AOI22XL U33633 ( .A0(n36107), .A1(n30366), .B0(n30358), .B1(n30392), .Y(
        n14757) );
  INVXL U33634 ( .A(filter_3[28]), .Y(n30367) );
  AOI22XL U33635 ( .A0(n36107), .A1(n30367), .B0(n30359), .B1(n30392), .Y(
        n14758) );
  INVXL U33636 ( .A(filter_3[29]), .Y(n30368) );
  AOI22XL U33637 ( .A0(n36107), .A1(n30368), .B0(n30360), .B1(n30392), .Y(
        n14759) );
  INVXL U33638 ( .A(filter_3[30]), .Y(n30369) );
  AOI22XL U33639 ( .A0(n36107), .A1(n30369), .B0(n30361), .B1(n30392), .Y(
        n14760) );
  INVXL U33640 ( .A(filter_3[31]), .Y(n30370) );
  AOI22XL U33641 ( .A0(n36107), .A1(n30370), .B0(n30362), .B1(n30392), .Y(
        n14761) );
  INVXL U33642 ( .A(filter_3[32]), .Y(n30371) );
  AOI22XL U33643 ( .A0(n36107), .A1(n30371), .B0(n30363), .B1(n30392), .Y(
        n14762) );
  AOI22XL U33644 ( .A0(n36107), .A1(n30365), .B0(n30364), .B1(n30392), .Y(
        n14749) );
  INVXL U33645 ( .A(filter_3[33]), .Y(n30372) );
  AOI22XL U33646 ( .A0(n36107), .A1(n30372), .B0(n30366), .B1(n30392), .Y(
        n14763) );
  INVXL U33647 ( .A(filter_3[34]), .Y(n30373) );
  AOI22XL U33648 ( .A0(n36107), .A1(n30373), .B0(n30367), .B1(n30392), .Y(
        n14764) );
  INVXL U33649 ( .A(filter_3[35]), .Y(n30374) );
  AOI22XL U33650 ( .A0(n36107), .A1(n30374), .B0(n30368), .B1(n30392), .Y(
        n14765) );
  INVXL U33651 ( .A(filter_3[36]), .Y(n30375) );
  AOI22XL U33652 ( .A0(n36107), .A1(n30375), .B0(n30369), .B1(n30392), .Y(
        n14766) );
  INVXL U33653 ( .A(filter_3[37]), .Y(n30376) );
  AOI22XL U33654 ( .A0(n36107), .A1(n30376), .B0(n30370), .B1(n30392), .Y(
        n14767) );
  INVXL U33655 ( .A(filter_3[38]), .Y(n30377) );
  AOI22XL U33656 ( .A0(n36107), .A1(n30377), .B0(n30371), .B1(n30392), .Y(
        n14768) );
  INVXL U33657 ( .A(filter_3[39]), .Y(n30379) );
  AOI22XL U33658 ( .A0(n36107), .A1(n30379), .B0(n30372), .B1(n30392), .Y(
        n14769) );
  INVXL U33659 ( .A(filter_3[40]), .Y(n30380) );
  AOI22XL U33660 ( .A0(n36107), .A1(n30380), .B0(n30373), .B1(n30392), .Y(
        n14770) );
  INVXL U33661 ( .A(filter_3[41]), .Y(n30381) );
  AOI22XL U33662 ( .A0(n36107), .A1(n30381), .B0(n30374), .B1(n30392), .Y(
        n14771) );
  INVXL U33663 ( .A(filter_3[42]), .Y(n30378) );
  AOI22XL U33664 ( .A0(n36107), .A1(n30378), .B0(n30375), .B1(n30392), .Y(
        n14772) );
  INVXL U33665 ( .A(filter_3[43]), .Y(n30383) );
  AOI22XL U33666 ( .A0(n36107), .A1(n30383), .B0(n30376), .B1(n30392), .Y(
        n14773) );
  INVXL U33667 ( .A(filter_3[44]), .Y(n30384) );
  AOI22XL U33668 ( .A0(n36107), .A1(n30384), .B0(n30377), .B1(n30392), .Y(
        n14774) );
  INVXL U33669 ( .A(filter_3[48]), .Y(n30390) );
  AOI22XL U33670 ( .A0(n36107), .A1(n30390), .B0(n30378), .B1(n30392), .Y(
        n14778) );
  INVXL U33671 ( .A(filter_3[45]), .Y(n30387) );
  AOI22XL U33672 ( .A0(n36107), .A1(n30387), .B0(n30379), .B1(n30392), .Y(
        n14775) );
  INVXL U33673 ( .A(filter_3[46]), .Y(n30388) );
  AOI22XL U33674 ( .A0(n36107), .A1(n30388), .B0(n30380), .B1(n30392), .Y(
        n14776) );
  INVXL U33675 ( .A(filter_3[47]), .Y(n30382) );
  AOI22XL U33676 ( .A0(n36107), .A1(n30382), .B0(n30381), .B1(n30392), .Y(
        n14777) );
  INVXL U33677 ( .A(filter_3[53]), .Y(n30391) );
  AOI22XL U33678 ( .A0(n36107), .A1(n30391), .B0(n30382), .B1(n30392), .Y(
        n14783) );
  INVXL U33679 ( .A(filter_3[50]), .Y(n30385) );
  AOI22XL U33680 ( .A0(n36107), .A1(n36142), .B0(n30385), .B1(n30392), .Y(
        n14786) );
  INVXL U33681 ( .A(filter_3[49]), .Y(n30386) );
  AOI22XL U33682 ( .A0(n36107), .A1(n30386), .B0(n30383), .B1(n30392), .Y(
        n14779) );
  AOI22XL U33683 ( .A0(n36107), .A1(n30385), .B0(n30384), .B1(n30392), .Y(
        n14780) );
  AOI22XL U33684 ( .A0(n36107), .A1(n36139), .B0(n30386), .B1(n30392), .Y(
        n14785) );
  INVXL U33685 ( .A(filter_3[51]), .Y(n30389) );
  AOI22XL U33686 ( .A0(n36107), .A1(n30389), .B0(n30387), .B1(n30392), .Y(
        n14781) );
  INVXL U33687 ( .A(filter_3[52]), .Y(n30393) );
  AOI22XL U33688 ( .A0(n36107), .A1(n30393), .B0(n30388), .B1(n30392), .Y(
        n14782) );
  AOI22XL U33689 ( .A0(n36107), .A1(n36145), .B0(n30389), .B1(n30392), .Y(
        n14787) );
  AOI22XL U33690 ( .A0(n36107), .A1(n36124), .B0(n30390), .B1(n30392), .Y(
        n14784) );
  AOI22XL U33691 ( .A0(n36107), .A1(n36151), .B0(n30391), .B1(n30392), .Y(
        n14789) );
  AOI22XL U33692 ( .A0(n36107), .A1(n36148), .B0(n30393), .B1(n30392), .Y(
        n14788) );
  INVXL U33693 ( .A(conv_2[437]), .Y(n30399) );
  NOR2BXL U33694 ( .AN(n30395), .B(n30394), .Y(n30397) );
  NAND2XL U33695 ( .A(conv_2[437]), .B(n30397), .Y(n30396) );
  OAI211XL U33696 ( .A0(conv_2[437]), .A1(n30397), .B0(n28751), .C0(n30396), 
        .Y(n30398) );
  OAI211XL U33697 ( .A0(n36070), .A1(n30399), .B0(n34621), .C0(n30398), .Y(
        n15282) );
  INVXL U33698 ( .A(conv_2[377]), .Y(n30405) );
  XOR2XL U33699 ( .A(n30401), .B(n30400), .Y(n30403) );
  NAND2XL U33700 ( .A(conv_2[377]), .B(n30403), .Y(n30402) );
  OAI211XL U33701 ( .A0(conv_2[377]), .A1(n30403), .B0(n33982), .C0(n30402), 
        .Y(n30404) );
  OAI211XL U33702 ( .A0(n36028), .A1(n30405), .B0(n34621), .C0(n30404), .Y(
        n15286) );
  INVXL U33703 ( .A(conv_2[17]), .Y(n30411) );
  XOR2XL U33704 ( .A(n30407), .B(n30406), .Y(n30409) );
  NAND2XL U33705 ( .A(conv_2[17]), .B(n30409), .Y(n30408) );
  OAI211XL U33706 ( .A0(conv_2[17]), .A1(n30409), .B0(n34028), .C0(n30408), 
        .Y(n30410) );
  OAI211XL U33707 ( .A0(n30412), .A1(n30411), .B0(n34621), .C0(n30410), .Y(
        n15310) );
  INVXL U33708 ( .A(conv_2[167]), .Y(n30416) );
  OAI211XL U33709 ( .A0(n30414), .A1(conv_2[167]), .B0(n31735), .C0(n30413), 
        .Y(n30415) );
  OAI211XL U33710 ( .A0(n34589), .A1(n30416), .B0(n34621), .C0(n30415), .Y(
        n15300) );
  INVXL U33711 ( .A(conv_2[77]), .Y(n30420) );
  OAI211XL U33712 ( .A0(n30418), .A1(conv_2[77]), .B0(n36020), .C0(n30417), 
        .Y(n30419) );
  OAI211XL U33713 ( .A0(n35879), .A1(n30420), .B0(n34621), .C0(n30419), .Y(
        n15306) );
  AOI22XL U33714 ( .A0(conv_2[538]), .A1(n30423), .B0(n30422), .B1(n30421), 
        .Y(n30425) );
  NAND2XL U33715 ( .A(conv_2[539]), .B(n30425), .Y(n30424) );
  OAI211XL U33716 ( .A0(conv_2[539]), .A1(n30425), .B0(n36020), .C0(n30424), 
        .Y(n30426) );
  OAI211XL U33717 ( .A0(n34789), .A1(n30427), .B0(n35859), .C0(n30426), .Y(
        n14844) );
  AOI2BB1XL U33718 ( .A0N(n33770), .A1N(n30435), .B0(n30436), .Y(n30432) );
  NAND2XL U33719 ( .A(conv_2[220]), .B(n30432), .Y(n30431) );
  OAI211XL U33720 ( .A0(conv_2[220]), .A1(n30432), .B0(n34028), .C0(n30431), 
        .Y(n30433) );
  OAI211XL U33721 ( .A0(n35934), .A1(n30434), .B0(n35859), .C0(n30433), .Y(
        n15058) );
  INVXL U33722 ( .A(conv_2[222]), .Y(n31122) );
  OAI21XL U33723 ( .A0(conv_2[220]), .A1(n30436), .B0(n33770), .Y(n35935) );
  AOI32XL U33724 ( .A0(conv_2[221]), .A1(n31121), .A2(n35936), .B0(n33770), 
        .B1(n35937), .Y(n30439) );
  NAND2XL U33725 ( .A(n31122), .B(n30439), .Y(n30438) );
  OAI211XL U33726 ( .A0(n31122), .A1(n30439), .B0(n34028), .C0(n30438), .Y(
        n30440) );
  OAI211XL U33727 ( .A0(n35934), .A1(n31122), .B0(n33815), .C0(n30440), .Y(
        n15056) );
  OAI32XL U33728 ( .A0(conv_2[133]), .A1(n30444), .A2(n30443), .B0(n30442), 
        .B1(n30441), .Y(n30446) );
  NAND2XL U33729 ( .A(conv_2[134]), .B(n30446), .Y(n30445) );
  OAI211XL U33730 ( .A0(conv_2[134]), .A1(n30446), .B0(n16657), .C0(n30445), 
        .Y(n30447) );
  OAI211XL U33731 ( .A0(n33853), .A1(n30448), .B0(n33815), .C0(n30447), .Y(
        n15114) );
  INVXL U33732 ( .A(conv_1[133]), .Y(n33041) );
  NAND4XL U33733 ( .A(conv_1[131]), .B(n30450), .C(conv_1[132]), .D(n30449), 
        .Y(n33043) );
  NAND2XL U33734 ( .A(n34292), .B(n30451), .Y(n33042) );
  NAND2XL U33735 ( .A(n33043), .B(n33042), .Y(n30453) );
  NAND2XL U33736 ( .A(conv_1[133]), .B(n30453), .Y(n30452) );
  OAI211XL U33737 ( .A0(conv_1[133]), .A1(n30453), .B0(n33822), .C0(n30452), 
        .Y(n30454) );
  OAI211XL U33738 ( .A0(n34296), .A1(n33041), .B0(n16652), .C0(n30454), .Y(
        n16330) );
  ADDFXL U33739 ( .A(conv_1[513]), .B(n30456), .CI(n30455), .CO(n27387), .S(
        n30457) );
  NAND2XL U33740 ( .A(n32656), .B(n30457), .Y(n30458) );
  OAI211XL U33741 ( .A0(n35547), .A1(n30459), .B0(n30458), .C0(n32867), .Y(
        n15950) );
  NAND2XL U33742 ( .A(conv_1[527]), .B(n30463), .Y(n30462) );
  OAI211XL U33743 ( .A0(conv_1[527]), .A1(n30463), .B0(n33788), .C0(n30462), 
        .Y(n30464) );
  OAI211XL U33744 ( .A0(n33432), .A1(n30465), .B0(n30464), .C0(n33542), .Y(
        n15936) );
  NAND2XL U33745 ( .A(conv_1[122]), .B(n30470), .Y(n30469) );
  OAI211XL U33746 ( .A0(conv_1[122]), .A1(n30470), .B0(n32181), .C0(n30469), 
        .Y(n30471) );
  OAI211XL U33747 ( .A0(n34296), .A1(n30472), .B0(n30471), .C0(n33542), .Y(
        n16341) );
  INVXL U33748 ( .A(conv_1[272]), .Y(n30478) );
  NAND2XL U33749 ( .A(conv_1[272]), .B(n30476), .Y(n30475) );
  OAI211XL U33750 ( .A0(conv_1[272]), .A1(n30476), .B0(n33982), .C0(n30475), 
        .Y(n30477) );
  OAI211XL U33751 ( .A0(n35426), .A1(n30478), .B0(n30477), .C0(n33542), .Y(
        n16191) );
  INVXL U33752 ( .A(conv_1[287]), .Y(n30484) );
  NAND2XL U33753 ( .A(conv_1[287]), .B(n30482), .Y(n30481) );
  OAI211XL U33754 ( .A0(conv_1[287]), .A1(n30482), .B0(n34028), .C0(n30481), 
        .Y(n30483) );
  OAI211XL U33755 ( .A0(n34325), .A1(n30484), .B0(n30483), .C0(n33542), .Y(
        n16176) );
  NAND2XL U33756 ( .A(conv_1[392]), .B(n30490), .Y(n30489) );
  OAI211XL U33757 ( .A0(conv_1[392]), .A1(n30490), .B0(n32181), .C0(n30489), 
        .Y(n30491) );
  OAI211XL U33758 ( .A0(n35477), .A1(n30492), .B0(n30491), .C0(n33542), .Y(
        n16071) );
  INVXL U33759 ( .A(conv_1[317]), .Y(n30496) );
  NAND2XL U33760 ( .A(conv_1[317]), .B(n30494), .Y(n30493) );
  OAI211XL U33761 ( .A0(conv_1[317]), .A1(n30494), .B0(n30090), .C0(n30493), 
        .Y(n30495) );
  OAI211XL U33762 ( .A0(n34263), .A1(n30496), .B0(n30495), .C0(n33542), .Y(
        n16146) );
  NOR2BXL U33763 ( .AN(n30498), .B(n30497), .Y(n30500) );
  NAND2XL U33764 ( .A(conv_3[482]), .B(n30500), .Y(n30499) );
  OAI211XL U33765 ( .A0(conv_3[482]), .A1(n30500), .B0(n32611), .C0(n30499), 
        .Y(n30501) );
  OAI211XL U33766 ( .A0(n35826), .A1(n30502), .B0(n30501), .C0(n35566), .Y(
        n15819) );
  INVXL U33767 ( .A(conv_3[527]), .Y(n30506) );
  NAND2XL U33768 ( .A(conv_3[527]), .B(n30504), .Y(n30503) );
  OAI211XL U33769 ( .A0(conv_3[527]), .A1(n30504), .B0(n36020), .C0(n30503), 
        .Y(n30505) );
  OAI211XL U33770 ( .A0(n31191), .A1(n30506), .B0(n30505), .C0(n35566), .Y(
        n15816) );
  INVXL U33771 ( .A(conv_3[452]), .Y(n30510) );
  NAND2XL U33772 ( .A(conv_3[452]), .B(n30508), .Y(n30507) );
  OAI211XL U33773 ( .A0(conv_3[452]), .A1(n30508), .B0(n31735), .C0(n30507), 
        .Y(n30509) );
  OAI211XL U33774 ( .A0(n35805), .A1(n30510), .B0(n30509), .C0(n35566), .Y(
        n15821) );
  NAND2XL U33775 ( .A(conv_3[347]), .B(n30515), .Y(n30514) );
  OAI211XL U33776 ( .A0(conv_3[347]), .A1(n30515), .B0(n24499), .C0(n30514), 
        .Y(n30516) );
  OAI211XL U33777 ( .A0(n34746), .A1(n30517), .B0(n30516), .C0(n35566), .Y(
        n15828) );
  INVXL U33778 ( .A(conv_3[511]), .Y(n30523) );
  AND2XL U33779 ( .A(n30519), .B(n30518), .Y(n30521) );
  NAND2XL U33780 ( .A(conv_3[511]), .B(n30521), .Y(n30520) );
  OAI211XL U33781 ( .A0(conv_3[511]), .A1(n30521), .B0(n32052), .C0(n30520), 
        .Y(n30522) );
  OAI211XL U33782 ( .A0(n33303), .A1(n30523), .B0(n30522), .C0(n33550), .Y(
        n15853) );
  NAND2XL U33783 ( .A(conv_3[481]), .B(n30527), .Y(n30526) );
  OAI211XL U33784 ( .A0(conv_3[481]), .A1(n30527), .B0(n33982), .C0(n30526), 
        .Y(n30528) );
  OAI211XL U33785 ( .A0(n35826), .A1(n30529), .B0(n30528), .C0(n33550), .Y(
        n15855) );
  INVXL U33786 ( .A(conv_3[211]), .Y(n30535) );
  NAND2XL U33787 ( .A(n30531), .B(n30530), .Y(n30533) );
  NAND2XL U33788 ( .A(n30535), .B(n30533), .Y(n30532) );
  OAI211XL U33789 ( .A0(n30535), .A1(n30533), .B0(n34028), .C0(n30532), .Y(
        n30534) );
  OAI211XL U33790 ( .A0(n35665), .A1(n30535), .B0(n30534), .C0(n33550), .Y(
        n15873) );
  NAND2XL U33791 ( .A(conv_3[286]), .B(n30540), .Y(n30539) );
  OAI211XL U33792 ( .A0(conv_3[286]), .A1(n30540), .B0(n33778), .C0(n30539), 
        .Y(n30541) );
  OAI211XL U33793 ( .A0(n35726), .A1(n30542), .B0(n30541), .C0(n33550), .Y(
        n15868) );
  NAND2XL U33794 ( .A(conv_3[407]), .B(n30546), .Y(n30545) );
  OAI211XL U33795 ( .A0(conv_3[407]), .A1(n30546), .B0(n16657), .C0(n30545), 
        .Y(n30547) );
  OAI211XL U33796 ( .A0(n34227), .A1(n30548), .B0(n30547), .C0(n35566), .Y(
        n15824) );
  NAND2XL U33797 ( .A(conv_3[17]), .B(n30553), .Y(n30552) );
  OAI211XL U33798 ( .A0(conv_3[17]), .A1(n30553), .B0(n32052), .C0(n30552), 
        .Y(n30554) );
  OAI211XL U33799 ( .A0(n35576), .A1(n30555), .B0(n30554), .C0(n35566), .Y(
        n15850) );
  INVXL U33800 ( .A(conv_3[316]), .Y(n30561) );
  NAND2XL U33801 ( .A(conv_3[316]), .B(n30559), .Y(n30558) );
  OAI211XL U33802 ( .A0(conv_3[316]), .A1(n30559), .B0(n33157), .C0(n30558), 
        .Y(n30560) );
  OAI211XL U33803 ( .A0(n35743), .A1(n30561), .B0(n30560), .C0(n33550), .Y(
        n15866) );
  INVXL U33804 ( .A(conv_3[361]), .Y(n30567) );
  NAND2XL U33805 ( .A(conv_3[361]), .B(n30565), .Y(n30564) );
  OAI211XL U33806 ( .A0(conv_3[361]), .A1(n30565), .B0(n33788), .C0(n30564), 
        .Y(n30566) );
  OAI211XL U33807 ( .A0(n35764), .A1(n30567), .B0(n30566), .C0(n33550), .Y(
        n15863) );
  INVXL U33808 ( .A(conv_3[346]), .Y(n30573) );
  NOR2BXL U33809 ( .AN(n30569), .B(n30568), .Y(n30571) );
  NAND2XL U33810 ( .A(conv_3[346]), .B(n30571), .Y(n30570) );
  OAI211XL U33811 ( .A0(conv_3[346]), .A1(n30571), .B0(n16656), .C0(n30570), 
        .Y(n30572) );
  OAI211XL U33812 ( .A0(n34746), .A1(n30573), .B0(n30572), .C0(n33550), .Y(
        n15864) );
  INVXL U33813 ( .A(conv_3[257]), .Y(n30579) );
  XOR2XL U33814 ( .A(n30575), .B(n30574), .Y(n30577) );
  NAND2XL U33815 ( .A(conv_3[257]), .B(n30577), .Y(n30576) );
  OAI211XL U33816 ( .A0(conv_3[257]), .A1(n30577), .B0(n34666), .C0(n30576), 
        .Y(n30578) );
  OAI211XL U33817 ( .A0(n35713), .A1(n30579), .B0(n30578), .C0(n35566), .Y(
        n15834) );
  INVXL U33818 ( .A(conv_1[437]), .Y(n30585) );
  XOR2XL U33819 ( .A(n30581), .B(n30580), .Y(n30583) );
  NAND2XL U33820 ( .A(conv_1[437]), .B(n30583), .Y(n30582) );
  OAI211XL U33821 ( .A0(conv_1[437]), .A1(n30583), .B0(n28751), .C0(n30582), 
        .Y(n30584) );
  OAI211XL U33822 ( .A0(n35520), .A1(n30585), .B0(n30584), .C0(n33542), .Y(
        n16026) );
  NOR2X1 U33823 ( .A(conv_1[27]), .B(n30589), .Y(n33203) );
  OAI21XL U33824 ( .A0(n33201), .A1(n33202), .B0(n30588), .Y(n30590) );
  AOI31XL U33825 ( .A0(n36020), .A1(n33203), .A2(n30590), .B0(n35549), .Y(
        n30593) );
  INVXL U33826 ( .A(n30589), .Y(n30591) );
  OAI2BB1XL U33827 ( .A0N(n30591), .A1N(n30590), .B0(n35336), .Y(n30592) );
  INVXL U33828 ( .A(conv_1[27]), .Y(n33200) );
  AOI32XL U33829 ( .A0(n35278), .A1(n30593), .A2(n30592), .B0(n33200), .B1(
        n30593), .Y(n16436) );
  OAI211XL U33830 ( .A0(n30595), .A1(conv_3[256]), .B0(n33778), .C0(n30594), 
        .Y(n30596) );
  OAI211XL U33831 ( .A0(n35713), .A1(n30597), .B0(n30596), .C0(n33550), .Y(
        n15870) );
  INVXL U33832 ( .A(conv_3[331]), .Y(n30601) );
  OAI211XL U33833 ( .A0(n30599), .A1(conv_3[331]), .B0(n16657), .C0(n30598), 
        .Y(n30600) );
  OAI211XL U33834 ( .A0(n35748), .A1(n30601), .B0(n30600), .C0(n33550), .Y(
        n15865) );
  OAI211XL U33835 ( .A0(conv_3[240]), .A1(n30603), .B0(n33788), .C0(n30602), 
        .Y(n30604) );
  OAI211XL U33836 ( .A0(n35706), .A1(n30605), .B0(n30604), .C0(n34755), .Y(
        n15907) );
  OAI211XL U33837 ( .A0(n30607), .A1(conv_3[255]), .B0(n27932), .C0(n30606), 
        .Y(n30608) );
  OAI211XL U33838 ( .A0(n35713), .A1(n30609), .B0(n30608), .C0(n34755), .Y(
        n15906) );
  INVXL U33839 ( .A(conv_3[315]), .Y(n30613) );
  OAI211XL U33840 ( .A0(n30611), .A1(conv_3[315]), .B0(n16656), .C0(n30610), 
        .Y(n30612) );
  OAI211XL U33841 ( .A0(n35743), .A1(n30613), .B0(n30612), .C0(n34755), .Y(
        n15902) );
  INVXL U33842 ( .A(conv_3[330]), .Y(n30617) );
  OAI211XL U33843 ( .A0(n30615), .A1(conv_3[330]), .B0(n32660), .C0(n30614), 
        .Y(n30616) );
  OAI211XL U33844 ( .A0(n35748), .A1(n30617), .B0(n30616), .C0(n34755), .Y(
        n15901) );
  INVXL U33845 ( .A(conv_3[285]), .Y(n30621) );
  OAI211XL U33846 ( .A0(conv_3[285]), .A1(n30619), .B0(n27932), .C0(n30618), 
        .Y(n30620) );
  OAI211XL U33847 ( .A0(n35726), .A1(n30621), .B0(n30620), .C0(n34755), .Y(
        n15904) );
  INVXL U33848 ( .A(conv_3[332]), .Y(n30627) );
  XOR2XL U33849 ( .A(n30623), .B(n30622), .Y(n30625) );
  NAND2XL U33850 ( .A(conv_3[332]), .B(n30625), .Y(n30624) );
  OAI211XL U33851 ( .A0(conv_3[332]), .A1(n30625), .B0(n32181), .C0(n30624), 
        .Y(n30626) );
  OAI211XL U33852 ( .A0(n35748), .A1(n30627), .B0(n30626), .C0(n35566), .Y(
        n15829) );
  INVXL U33853 ( .A(conv_3[212]), .Y(n30631) );
  NAND2XL U33854 ( .A(conv_3[212]), .B(n30629), .Y(n30628) );
  OAI211XL U33855 ( .A0(conv_3[212]), .A1(n30629), .B0(n33712), .C0(n30628), 
        .Y(n30630) );
  OAI211XL U33856 ( .A0(n35665), .A1(n30631), .B0(n30630), .C0(n35566), .Y(
        n15837) );
  INVXL U33857 ( .A(conv_3[406]), .Y(n30635) );
  OAI211XL U33858 ( .A0(conv_3[406]), .A1(n30633), .B0(n34666), .C0(n30632), 
        .Y(n30634) );
  OAI211XL U33859 ( .A0(n34227), .A1(n30635), .B0(n30634), .C0(n33550), .Y(
        n15860) );
  INVXL U33860 ( .A(conv_3[376]), .Y(n30639) );
  NAND2XL U33861 ( .A(conv_3[376]), .B(n30637), .Y(n30636) );
  OAI211XL U33862 ( .A0(conv_3[376]), .A1(n30637), .B0(n33822), .C0(n30636), 
        .Y(n30638) );
  OAI211XL U33863 ( .A0(n34168), .A1(n30639), .B0(n30638), .C0(n33550), .Y(
        n15862) );
  INVXL U33864 ( .A(conv_3[271]), .Y(n30643) );
  NAND2XL U33865 ( .A(conv_3[271]), .B(n30641), .Y(n30640) );
  OAI211XL U33866 ( .A0(conv_3[271]), .A1(n30641), .B0(n16656), .C0(n30640), 
        .Y(n30642) );
  OAI211XL U33867 ( .A0(n34709), .A1(n30643), .B0(n30642), .C0(n33550), .Y(
        n15869) );
  AOI22XL U33868 ( .A0(n34821), .A1(n30645), .B0(n30644), .B1(n34817), .Y(
        N29244) );
  AOI22XL U33869 ( .A0(n34821), .A1(n30647), .B0(n30646), .B1(n34817), .Y(
        N29245) );
  OAI211XL U33870 ( .A0(conv_1[390]), .A1(n30649), .B0(n33822), .C0(n30648), 
        .Y(n30650) );
  OAI211XL U33871 ( .A0(n35477), .A1(n30651), .B0(n30650), .C0(n34773), .Y(
        n16073) );
  INVXL U33872 ( .A(conv_1[270]), .Y(n30655) );
  OAI211XL U33873 ( .A0(conv_1[270]), .A1(n30653), .B0(n34666), .C0(n30652), 
        .Y(n30654) );
  OAI211XL U33874 ( .A0(n35426), .A1(n30655), .B0(n30654), .C0(n34773), .Y(
        n16193) );
  INVXL U33875 ( .A(conv_1[436]), .Y(n30661) );
  NAND2XL U33876 ( .A(n30657), .B(n30656), .Y(n30659) );
  NAND2XL U33877 ( .A(n30661), .B(n30659), .Y(n30658) );
  OAI211XL U33878 ( .A0(n30661), .A1(n30659), .B0(n33822), .C0(n30658), .Y(
        n30660) );
  OAI211XL U33879 ( .A0(n35520), .A1(n30661), .B0(n30660), .C0(n33067), .Y(
        n16027) );
  INVXL U33880 ( .A(conv_1[435]), .Y(n30665) );
  OAI211XL U33881 ( .A0(n30663), .A1(conv_1[435]), .B0(n33822), .C0(n30662), 
        .Y(n30664) );
  OAI211XL U33882 ( .A0(n35520), .A1(n30665), .B0(n30664), .C0(n34773), .Y(
        n16028) );
  NOR2BXL U33883 ( .AN(n30667), .B(n30666), .Y(n30669) );
  NAND2XL U33884 ( .A(conv_1[391]), .B(n30669), .Y(n30668) );
  OAI211XL U33885 ( .A0(conv_1[391]), .A1(n30669), .B0(n28751), .C0(n30668), 
        .Y(n30670) );
  OAI211XL U33886 ( .A0(n35477), .A1(n30671), .B0(n30670), .C0(n33067), .Y(
        n16072) );
  INVXL U33887 ( .A(conv_1[421]), .Y(n33399) );
  NAND2XL U33888 ( .A(n30672), .B(conv_1[420]), .Y(n30673) );
  OAI2BB1XL U33889 ( .A0N(n35272), .A1N(n30673), .B0(n34768), .Y(n33398) );
  OR2XL U33890 ( .A(n30673), .B(n35499), .Y(n34770) );
  NAND2XL U33891 ( .A(conv_1[421]), .B(n30675), .Y(n30674) );
  OAI211XL U33892 ( .A0(conv_1[421]), .A1(n30675), .B0(n32181), .C0(n30674), 
        .Y(n30676) );
  OAI211XL U33893 ( .A0(n35504), .A1(n33399), .B0(n30676), .C0(n33067), .Y(
        n16042) );
  INVXL U33894 ( .A(conv_1[271]), .Y(n30680) );
  OAI211XL U33895 ( .A0(conv_1[271]), .A1(n30678), .B0(n32181), .C0(n30677), 
        .Y(n30679) );
  OAI211XL U33896 ( .A0(n35426), .A1(n30680), .B0(n30679), .C0(n33067), .Y(
        n16192) );
  INVXL U33897 ( .A(conv_1[526]), .Y(n30684) );
  OAI211XL U33898 ( .A0(conv_1[526]), .A1(n30682), .B0(n33778), .C0(n30681), 
        .Y(n30683) );
  OAI211XL U33899 ( .A0(n33432), .A1(n30684), .B0(n30683), .C0(n33067), .Y(
        n15937) );
  INVXL U33900 ( .A(conv_1[286]), .Y(n30688) );
  OAI211XL U33901 ( .A0(conv_1[286]), .A1(n30686), .B0(n33982), .C0(n30685), 
        .Y(n30687) );
  OAI211XL U33902 ( .A0(n34325), .A1(n30688), .B0(n30687), .C0(n33067), .Y(
        n16177) );
  AOI21XL U33903 ( .A0(n33878), .A1(n30690), .B0(n30689), .Y(n30692) );
  NAND2XL U33904 ( .A(conv_3[234]), .B(n30692), .Y(n30691) );
  OAI211XL U33905 ( .A0(conv_3[234]), .A1(n30692), .B0(n33912), .C0(n30691), 
        .Y(n30693) );
  OAI211XL U33906 ( .A0(n35676), .A1(n30694), .B0(n16649), .C0(n30693), .Y(
        n15589) );
  NAND2XL U33907 ( .A(conv_1[499]), .B(n30698), .Y(n30697) );
  OAI211XL U33908 ( .A0(conv_1[499]), .A1(n30698), .B0(n34666), .C0(n30697), 
        .Y(n30699) );
  OAI211XL U33909 ( .A0(n33427), .A1(n30700), .B0(n35489), .C0(n30699), .Y(
        n15964) );
  INVXL U33910 ( .A(conv_3[32]), .Y(n30706) );
  NAND2XL U33911 ( .A(n30702), .B(n30701), .Y(n30704) );
  NAND2XL U33912 ( .A(n30706), .B(n30704), .Y(n30703) );
  OAI211XL U33913 ( .A0(n30706), .A1(n30704), .B0(n27932), .C0(n30703), .Y(
        n30705) );
  OAI211XL U33914 ( .A0(n35594), .A1(n30706), .B0(n35566), .C0(n30705), .Y(
        n15849) );
  INVXL U33915 ( .A(conv_3[137]), .Y(n30712) );
  NAND2XL U33916 ( .A(n30708), .B(n30707), .Y(n30710) );
  NAND2XL U33917 ( .A(n30712), .B(n30710), .Y(n30709) );
  OAI211XL U33918 ( .A0(n30712), .A1(n30710), .B0(n36020), .C0(n30709), .Y(
        n30711) );
  OAI211XL U33919 ( .A0(n34737), .A1(n30712), .B0(n35566), .C0(n30711), .Y(
        n15842) );
  INVXL U33920 ( .A(conv_3[302]), .Y(n30718) );
  NAND2XL U33921 ( .A(n30714), .B(n30713), .Y(n30716) );
  NAND2XL U33922 ( .A(n30718), .B(n30716), .Y(n30715) );
  OAI211XL U33923 ( .A0(n30718), .A1(n30716), .B0(n32660), .C0(n30715), .Y(
        n30717) );
  OAI211XL U33924 ( .A0(n35736), .A1(n30718), .B0(n35566), .C0(n30717), .Y(
        n15831) );
  INVXL U33925 ( .A(conv_3[512]), .Y(n30722) );
  NAND2XL U33926 ( .A(conv_3[512]), .B(n30720), .Y(n30719) );
  OAI211XL U33927 ( .A0(conv_3[512]), .A1(n30720), .B0(n27932), .C0(n30719), 
        .Y(n30721) );
  OAI211XL U33928 ( .A0(n33303), .A1(n30722), .B0(n35566), .C0(n30721), .Y(
        n15817) );
  INVXL U33929 ( .A(conv_3[497]), .Y(n30728) );
  NOR2BXL U33930 ( .AN(n30724), .B(n30723), .Y(n30726) );
  NAND2XL U33931 ( .A(conv_3[497]), .B(n30726), .Y(n30725) );
  OAI211XL U33932 ( .A0(conv_3[497]), .A1(n30726), .B0(n34666), .C0(n30725), 
        .Y(n30727) );
  OAI211XL U33933 ( .A0(n35841), .A1(n30728), .B0(n35566), .C0(n30727), .Y(
        n15818) );
  INVXL U33934 ( .A(conv_3[496]), .Y(n30734) );
  NOR2BXL U33935 ( .AN(n30730), .B(n30729), .Y(n30732) );
  NAND2XL U33936 ( .A(conv_3[496]), .B(n30732), .Y(n30731) );
  OAI211XL U33937 ( .A0(conv_3[496]), .A1(n30732), .B0(n16656), .C0(n30731), 
        .Y(n30733) );
  OAI211XL U33938 ( .A0(n35841), .A1(n30734), .B0(n33550), .C0(n30733), .Y(
        n15854) );
  INVXL U33939 ( .A(conv_1[407]), .Y(n30740) );
  XOR2XL U33940 ( .A(n30736), .B(n30735), .Y(n30738) );
  NAND2XL U33941 ( .A(conv_1[407]), .B(n30738), .Y(n30737) );
  OAI211XL U33942 ( .A0(conv_1[407]), .A1(n30738), .B0(n35336), .C0(n30737), 
        .Y(n30739) );
  OAI211XL U33943 ( .A0(n35487), .A1(n30740), .B0(n33542), .C0(n30739), .Y(
        n16056) );
  INVXL U33944 ( .A(conv_3[122]), .Y(n30746) );
  NAND2XL U33945 ( .A(conv_3[122]), .B(n30744), .Y(n30743) );
  OAI211XL U33946 ( .A0(conv_3[122]), .A1(n30744), .B0(n34666), .C0(n30743), 
        .Y(n30745) );
  OAI211XL U33947 ( .A0(n35626), .A1(n30746), .B0(n35566), .C0(n30745), .Y(
        n15843) );
  INVXL U33948 ( .A(conv_3[47]), .Y(n30752) );
  NAND2XL U33949 ( .A(conv_3[47]), .B(n30750), .Y(n30749) );
  OAI211XL U33950 ( .A0(conv_3[47]), .A1(n30750), .B0(n32611), .C0(n30749), 
        .Y(n30751) );
  OAI211XL U33951 ( .A0(n34392), .A1(n30752), .B0(n35566), .C0(n30751), .Y(
        n15848) );
  INVXL U33952 ( .A(conv_1[124]), .Y(n30758) );
  NAND2XL U33953 ( .A(conv_1[124]), .B(n30756), .Y(n30755) );
  OAI211XL U33954 ( .A0(conv_1[124]), .A1(n30756), .B0(n32181), .C0(n30755), 
        .Y(n30757) );
  OAI211XL U33955 ( .A0(n34296), .A1(n30758), .B0(n35489), .C0(n30757), .Y(
        n16339) );
  NAND2XL U33956 ( .A(conv_1[394]), .B(n30762), .Y(n30761) );
  OAI211XL U33957 ( .A0(conv_1[394]), .A1(n30762), .B0(n33822), .C0(n30761), 
        .Y(n30763) );
  OAI211XL U33958 ( .A0(n35477), .A1(n30764), .B0(n35489), .C0(n30763), .Y(
        n16069) );
  AOI21XL U33959 ( .A0(n30767), .A1(n30766), .B0(n30765), .Y(n30769) );
  NAND2XL U33960 ( .A(conv_1[274]), .B(n30769), .Y(n30768) );
  OAI211XL U33961 ( .A0(conv_1[274]), .A1(n30769), .B0(n31735), .C0(n30768), 
        .Y(n30770) );
  OAI211XL U33962 ( .A0(n35426), .A1(n30771), .B0(n35489), .C0(n30770), .Y(
        n16189) );
  AOI21XL U33963 ( .A0(n30774), .A1(n30773), .B0(n30772), .Y(n30776) );
  NAND2XL U33964 ( .A(conv_1[289]), .B(n30776), .Y(n30775) );
  OAI211XL U33965 ( .A0(conv_1[289]), .A1(n30776), .B0(n32660), .C0(n30775), 
        .Y(n30777) );
  OAI211XL U33966 ( .A0(n34325), .A1(n30778), .B0(n35489), .C0(n30777), .Y(
        n16174) );
  INVXL U33967 ( .A(conv_3[467]), .Y(n30784) );
  XOR2XL U33968 ( .A(n30780), .B(n30779), .Y(n30782) );
  NAND2XL U33969 ( .A(conv_3[467]), .B(n30782), .Y(n30781) );
  OAI211XL U33970 ( .A0(conv_3[467]), .A1(n30782), .B0(n33982), .C0(n30781), 
        .Y(n30783) );
  OAI211XL U33971 ( .A0(n35813), .A1(n30784), .B0(n35566), .C0(n30783), .Y(
        n15820) );
  INVXL U33972 ( .A(conv_3[2]), .Y(n30788) );
  NAND2XL U33973 ( .A(conv_3[2]), .B(n30786), .Y(n30785) );
  OAI211XL U33974 ( .A0(conv_3[2]), .A1(n30786), .B0(n33778), .C0(n30785), .Y(
        n30787) );
  OAI211XL U33975 ( .A0(n34383), .A1(n30788), .B0(n35566), .C0(n30787), .Y(
        n15851) );
  OAI211XL U33976 ( .A0(n30790), .A1(conv_3[466]), .B0(n31735), .C0(n30789), 
        .Y(n30791) );
  OAI211XL U33977 ( .A0(n35813), .A1(n30792), .B0(n33550), .C0(n30791), .Y(
        n15856) );
  INVXL U33978 ( .A(conv_3[107]), .Y(n30798) );
  XOR2XL U33979 ( .A(n30794), .B(n30793), .Y(n30796) );
  NAND2XL U33980 ( .A(conv_3[107]), .B(n30796), .Y(n30795) );
  OAI211XL U33981 ( .A0(conv_3[107]), .A1(n30796), .B0(n33712), .C0(n30795), 
        .Y(n30797) );
  OAI211XL U33982 ( .A0(n34200), .A1(n30798), .B0(n35566), .C0(n30797), .Y(
        n15844) );
  INVXL U33983 ( .A(conv_3[197]), .Y(n30804) );
  XOR2XL U33984 ( .A(n30800), .B(n30799), .Y(n30802) );
  NAND2XL U33985 ( .A(conv_3[197]), .B(n30802), .Y(n30801) );
  OAI211XL U33986 ( .A0(conv_3[197]), .A1(n30802), .B0(n27932), .C0(n30801), 
        .Y(n30803) );
  OAI211XL U33987 ( .A0(n35646), .A1(n30804), .B0(n35566), .C0(n30803), .Y(
        n15838) );
  NAND2XL U33988 ( .A(conv_3[422]), .B(n30808), .Y(n30807) );
  OAI211XL U33989 ( .A0(conv_3[422]), .A1(n30808), .B0(n16657), .C0(n30807), 
        .Y(n30809) );
  OAI211XL U33990 ( .A0(n35778), .A1(n30810), .B0(n35566), .C0(n30809), .Y(
        n15823) );
  XOR2XL U33991 ( .A(n30812), .B(n30811), .Y(n30814) );
  NAND2XL U33992 ( .A(conv_3[437]), .B(n30814), .Y(n30813) );
  OAI211XL U33993 ( .A0(conv_3[437]), .A1(n30814), .B0(n33982), .C0(n30813), 
        .Y(n30815) );
  OAI211XL U33994 ( .A0(n35792), .A1(n30816), .B0(n35566), .C0(n30815), .Y(
        n15822) );
  INVXL U33995 ( .A(conv_3[152]), .Y(n30822) );
  XOR2XL U33996 ( .A(n30818), .B(n30817), .Y(n30820) );
  NAND2XL U33997 ( .A(conv_3[152]), .B(n30820), .Y(n30819) );
  OAI211XL U33998 ( .A0(conv_3[152]), .A1(n30820), .B0(n27932), .C0(n30819), 
        .Y(n30821) );
  OAI211XL U33999 ( .A0(n34751), .A1(n30822), .B0(n35566), .C0(n30821), .Y(
        n15841) );
  INVXL U34000 ( .A(conv_3[92]), .Y(n30828) );
  XOR2XL U34001 ( .A(n30824), .B(n30823), .Y(n30826) );
  NAND2XL U34002 ( .A(conv_3[92]), .B(n30826), .Y(n30825) );
  OAI211XL U34003 ( .A0(conv_3[92]), .A1(n30826), .B0(n34028), .C0(n30825), 
        .Y(n30827) );
  OAI211XL U34004 ( .A0(n35618), .A1(n30828), .B0(n35566), .C0(n30827), .Y(
        n15845) );
  OAI211XL U34005 ( .A0(n30830), .A1(conv_3[105]), .B0(n33778), .C0(n30829), 
        .Y(n30831) );
  OAI211XL U34006 ( .A0(n34200), .A1(n30832), .B0(n34755), .C0(n30831), .Y(
        n15916) );
  OAI211XL U34007 ( .A0(n30834), .A1(conv_3[90]), .B0(n34666), .C0(n30833), 
        .Y(n30835) );
  OAI211XL U34008 ( .A0(n35618), .A1(n30836), .B0(n34755), .C0(n30835), .Y(
        n15917) );
  INVXL U34009 ( .A(conv_3[120]), .Y(n30840) );
  OAI211XL U34010 ( .A0(n30838), .A1(conv_3[120]), .B0(n34666), .C0(n30837), 
        .Y(n30839) );
  OAI211XL U34011 ( .A0(n35626), .A1(n30840), .B0(n34755), .C0(n30839), .Y(
        n15915) );
  INVXL U34012 ( .A(conv_3[195]), .Y(n30844) );
  OAI211XL U34013 ( .A0(n30842), .A1(conv_3[195]), .B0(n27932), .C0(n30841), 
        .Y(n30843) );
  OAI211XL U34014 ( .A0(n35646), .A1(n30844), .B0(n34755), .C0(n30843), .Y(
        n15910) );
  XOR2XL U34015 ( .A(n30846), .B(n30845), .Y(n30848) );
  NAND2XL U34016 ( .A(conv_3[227]), .B(n30848), .Y(n30847) );
  OAI211XL U34017 ( .A0(conv_3[227]), .A1(n30848), .B0(n27932), .C0(n30847), 
        .Y(n30849) );
  OAI211XL U34018 ( .A0(n35676), .A1(n30850), .B0(n35566), .C0(n30849), .Y(
        n15836) );
  INVXL U34019 ( .A(conv_3[392]), .Y(n30856) );
  XOR2XL U34020 ( .A(n30852), .B(n30851), .Y(n30854) );
  NAND2XL U34021 ( .A(conv_3[392]), .B(n30854), .Y(n30853) );
  OAI211XL U34022 ( .A0(conv_3[392]), .A1(n30854), .B0(n33778), .C0(n30853), 
        .Y(n30855) );
  OAI211XL U34023 ( .A0(n33703), .A1(n30856), .B0(n35566), .C0(n30855), .Y(
        n15825) );
  OAI21XL U34024 ( .A0(n30860), .A1(n36042), .B0(n35976), .Y(n30859) );
  NAND2XL U34025 ( .A(n30862), .B(n34735), .Y(n15003) );
  ADDFX1 U34026 ( .A(conv_2[488]), .B(n34132), .CI(n30863), .CO(n27753), .S(
        n30864) );
  AOI22XL U34027 ( .A0(n16656), .A1(n30864), .B0(conv_2[488]), .B1(n33598), 
        .Y(n30865) );
  NAND2XL U34028 ( .A(n30865), .B(n34735), .Y(n14880) );
  NAND2XL U34029 ( .A(n30866), .B(n30961), .Y(n30868) );
  AOI211XL U34030 ( .A0(n30870), .A1(n30868), .B0(n36042), .C0(n30867), .Y(
        n30869) );
  AOI2BB1XL U34031 ( .A0N(n30870), .A1N(n36070), .B0(n30869), .Y(n30871) );
  NAND2XL U34032 ( .A(n30871), .B(n34735), .Y(n14907) );
  ADDFXL U34033 ( .A(conv_2[52]), .B(n31137), .CI(n30872), .CO(n27814), .S(
        n30874) );
  AOI22XL U34034 ( .A0(n32611), .A1(n30874), .B0(conv_2[52]), .B1(n30873), .Y(
        n30875) );
  NAND2XL U34035 ( .A(n30875), .B(n34735), .Y(n15171) );
  AOI32XL U34036 ( .A0(conv_2[455]), .A1(n30877), .A2(n30876), .B0(n33611), 
        .B1(n30877), .Y(n30879) );
  AOI211XL U34037 ( .A0(n30881), .A1(n30879), .B0(n36042), .C0(n30878), .Y(
        n30880) );
  AOI2BB1XL U34038 ( .A0N(n30881), .A1N(n34441), .B0(n30880), .Y(n30882) );
  NAND2XL U34039 ( .A(n30882), .B(n34735), .Y(n14902) );
  AOI21XL U34040 ( .A0(n33691), .A1(conv_2[414]), .B0(n36045), .Y(n36038) );
  AOI22XL U34041 ( .A0(n33778), .A1(n30886), .B0(conv_2[416]), .B1(n33687), 
        .Y(n30887) );
  NAND2XL U34042 ( .A(n30887), .B(n34735), .Y(n14927) );
  OAI21XL U34043 ( .A0(n30891), .A1(n36042), .B0(n35963), .Y(n30890) );
  NAND2XL U34044 ( .A(n30893), .B(n34735), .Y(n15013) );
  NAND2XL U34045 ( .A(n29831), .B(n30894), .Y(n30896) );
  AOI21X1 U34046 ( .A0(n30897), .A1(n30896), .B0(n30895), .Y(n33973) );
  AOI22XL U34047 ( .A0(n33982), .A1(n30898), .B0(conv_2[176]), .B1(n30969), 
        .Y(n30899) );
  NAND2XL U34048 ( .A(n30899), .B(n34735), .Y(n15087) );
  OAI21XL U34049 ( .A0(n30903), .A1(n16655), .B0(n34177), .Y(n30902) );
  AOI32XL U34050 ( .A0(n36020), .A1(n30904), .A2(n30903), .B0(conv_2[474]), 
        .B1(n30902), .Y(n30905) );
  NAND2XL U34051 ( .A(n30905), .B(n34735), .Y(n14889) );
  ADDFX1 U34052 ( .A(conv_2[174]), .B(n29831), .CI(n30906), .CO(n30894), .S(
        n30907) );
  AOI22XL U34053 ( .A0(n34028), .A1(n30907), .B0(conv_2[174]), .B1(n30969), 
        .Y(n30908) );
  NAND2XL U34054 ( .A(n30908), .B(n34735), .Y(n15089) );
  INVXL U34055 ( .A(conv_2[506]), .Y(n33168) );
  OAI21XL U34056 ( .A0(conv_2[505]), .A1(n36086), .B0(n36088), .Y(n33167) );
  INVXL U34057 ( .A(conv_2[504]), .Y(n36083) );
  NAND2XL U34058 ( .A(conv_2[503]), .B(n36074), .Y(n36080) );
  OAI2BB1XL U34059 ( .A0N(conv_2[505]), .A1N(n36087), .B0(n36081), .Y(n33704)
         );
  NAND2XL U34060 ( .A(n33167), .B(n33704), .Y(n30913) );
  AOI211XL U34061 ( .A0(n33168), .A1(n30913), .B0(n36042), .C0(n30912), .Y(
        n30914) );
  AOI2BB1XL U34062 ( .A0N(n33168), .A1N(n36091), .B0(n30914), .Y(n30915) );
  NAND2XL U34063 ( .A(n30915), .B(n34735), .Y(n14867) );
  INVXL U34064 ( .A(conv_2[294]), .Y(n30922) );
  NAND2XL U34065 ( .A(n35957), .B(n30979), .Y(n30918) );
  OAI21XL U34066 ( .A0(n35957), .A1(n30979), .B0(n30918), .Y(n30920) );
  AOI211XL U34067 ( .A0(n30922), .A1(n30920), .B0(n16655), .C0(n30919), .Y(
        n30921) );
  AOI2BB1XL U34068 ( .A0N(n30922), .A1N(n35963), .B0(n30921), .Y(n30923) );
  NAND2XL U34069 ( .A(n30923), .B(n34735), .Y(n15009) );
  INVXL U34070 ( .A(conv_2[88]), .Y(n32671) );
  NAND3XL U34071 ( .A(n30925), .B(conv_2[87]), .C(n30924), .Y(n32673) );
  NAND3XL U34072 ( .A(n30927), .B(n35876), .C(n30926), .Y(n32672) );
  OAI21XL U34073 ( .A0(n16654), .A1(n30929), .B0(n35879), .Y(n30928) );
  NAND2XL U34074 ( .A(n30930), .B(n34735), .Y(n15145) );
  NAND2BXL U34075 ( .AN(n30932), .B(n30931), .Y(n30934) );
  AOI211XL U34076 ( .A0(n30936), .A1(n30934), .B0(n36042), .C0(n30933), .Y(
        n30935) );
  AOI2BB1XL U34077 ( .A0N(n30936), .A1N(n34458), .B0(n30935), .Y(n30937) );
  NAND2XL U34078 ( .A(n30937), .B(n34735), .Y(n15047) );
  OAI2BB1XL U34079 ( .A0N(n30940), .A1N(n30939), .B0(n30938), .Y(n30942) );
  AOI211XL U34080 ( .A0(n30944), .A1(n30942), .B0(n16654), .C0(n30941), .Y(
        n30943) );
  AOI2BB1XL U34081 ( .A0N(n30944), .A1N(n34447), .B0(n30943), .Y(n30945) );
  NAND2XL U34082 ( .A(n30945), .B(n34735), .Y(n15139) );
  AOI22XL U34083 ( .A0(n35914), .A1(n30948), .B0(n30947), .B1(n30946), .Y(
        n30950) );
  AOI211XL U34084 ( .A0(n30952), .A1(n30950), .B0(n36042), .C0(n30949), .Y(
        n30951) );
  NAND2XL U34085 ( .A(n30953), .B(n34735), .Y(n15076) );
  OAI21XL U34086 ( .A0(n33571), .A1(intadd_0_n1), .B0(n30954), .Y(n30956) );
  AOI211XL U34087 ( .A0(n30959), .A1(n30956), .B0(n36001), .C0(n30955), .Y(
        n30957) );
  AOI2BB1XL U34088 ( .A0N(n30959), .A1N(n30958), .B0(n30957), .Y(n30960) );
  NAND2XL U34089 ( .A(n30960), .B(n34735), .Y(n15203) );
  AOI32XL U34090 ( .A0(conv_2[446]), .A1(n30962), .A2(n30961), .B0(n36067), 
        .B1(n30962), .Y(n30964) );
  AOI211XL U34091 ( .A0(n30966), .A1(n30964), .B0(n36042), .C0(n30963), .Y(
        n30965) );
  AOI2BB1XL U34092 ( .A0N(n30966), .A1N(n36070), .B0(n30965), .Y(n30967) );
  NAND2XL U34093 ( .A(n30967), .B(n34735), .Y(n14906) );
  AOI22XL U34094 ( .A0(n32052), .A1(n30970), .B0(conv_2[171]), .B1(n30969), 
        .Y(n30971) );
  NAND2XL U34095 ( .A(n30971), .B(n34735), .Y(n15092) );
  OAI21XL U34096 ( .A0(n33735), .A1(n30973), .B0(n30972), .Y(n30975) );
  AOI211XL U34097 ( .A0(n30977), .A1(n30975), .B0(n36001), .C0(n30974), .Y(
        n30976) );
  AOI2BB1XL U34098 ( .A0N(n30977), .A1N(n35846), .B0(n30976), .Y(n30978) );
  NAND2XL U34099 ( .A(n30978), .B(n34735), .Y(n15159) );
  OAI21XL U34100 ( .A0(conv_2[294]), .A1(n30979), .B0(n35957), .Y(n35962) );
  AOI22XL U34101 ( .A0(n32656), .A1(n30980), .B0(conv_2[296]), .B1(n35959), 
        .Y(n30981) );
  NAND2XL U34102 ( .A(n30981), .B(n34735), .Y(n15007) );
  ADDFXL U34103 ( .A(conv_2[530]), .B(n33629), .CI(n30982), .CO(n29625), .S(
        n30983) );
  AOI22XL U34104 ( .A0(n34028), .A1(n30983), .B0(conv_2[530]), .B1(n33624), 
        .Y(n30984) );
  NAND2XL U34105 ( .A(n30984), .B(n34735), .Y(n14853) );
  AOI32XL U34106 ( .A0(conv_2[281]), .A1(n30986), .A2(n30985), .B0(n35950), 
        .B1(n30986), .Y(n30988) );
  AOI211XL U34107 ( .A0(n30990), .A1(n30988), .B0(n36042), .C0(n30987), .Y(
        n30989) );
  AOI2BB1XL U34108 ( .A0N(n30990), .A1N(n30994), .B0(n30989), .Y(n30991) );
  NAND2XL U34109 ( .A(n30991), .B(n34735), .Y(n15016) );
  NAND2XL U34110 ( .A(n30993), .B(n30992), .Y(n30996) );
  OAI21XL U34111 ( .A0(n16654), .A1(n30996), .B0(n30994), .Y(n30995) );
  NAND2XL U34112 ( .A(n30998), .B(n34735), .Y(n15015) );
  ADDFX1 U34113 ( .A(conv_2[293]), .B(n35957), .CI(n30999), .CO(n30979), .S(
        n31000) );
  AOI22XL U34114 ( .A0(n36056), .A1(n31000), .B0(conv_2[293]), .B1(n35959), 
        .Y(n31001) );
  NAND2XL U34115 ( .A(n31001), .B(n34735), .Y(n15010) );
  INVXL U34116 ( .A(conv_2[86]), .Y(n31006) );
  OAI21XL U34117 ( .A0(n31005), .A1(n16655), .B0(n35879), .Y(n31004) );
  AOI32XL U34118 ( .A0(n31735), .A1(n31006), .A2(n31005), .B0(conv_2[86]), 
        .B1(n31004), .Y(n31007) );
  NAND2XL U34119 ( .A(n31007), .B(n34735), .Y(n15147) );
  NAND2XL U34120 ( .A(n31009), .B(n31008), .Y(n31011) );
  AOI211XL U34121 ( .A0(n31014), .A1(n31011), .B0(n36042), .C0(n31010), .Y(
        n31012) );
  NAND2XL U34122 ( .A(n31015), .B(n34735), .Y(n14857) );
  INVXL U34123 ( .A(conv_2[500]), .Y(n31020) );
  OAI21XL U34124 ( .A0(n31019), .A1(n16654), .B0(n36091), .Y(n31018) );
  AOI32XL U34125 ( .A0(n24378), .A1(n31020), .A2(n31019), .B0(conv_2[500]), 
        .B1(n31018), .Y(n31021) );
  NAND2XL U34126 ( .A(n31021), .B(n34735), .Y(n14873) );
  INVXL U34127 ( .A(conv_3[301]), .Y(n31025) );
  OAI211XL U34128 ( .A0(n31023), .A1(conv_3[301]), .B0(n32181), .C0(n31022), 
        .Y(n31024) );
  OAI211XL U34129 ( .A0(n35736), .A1(n31025), .B0(n33550), .C0(n31024), .Y(
        n15867) );
  INVXL U34130 ( .A(conv_3[0]), .Y(n31029) );
  OAI211XL U34131 ( .A0(conv_3[0]), .A1(n31027), .B0(n27932), .C0(n31026), .Y(
        n31028) );
  OAI211XL U34132 ( .A0(n34383), .A1(n31029), .B0(n34755), .C0(n31028), .Y(
        n15923) );
  OAI211XL U34133 ( .A0(n31031), .A1(conv_3[436]), .B0(n33778), .C0(n31030), 
        .Y(n31032) );
  OAI211XL U34134 ( .A0(n35792), .A1(n31033), .B0(n33550), .C0(n31032), .Y(
        n15858) );
  INVXL U34135 ( .A(conv_3[391]), .Y(n31037) );
  OAI211XL U34136 ( .A0(n31035), .A1(conv_3[391]), .B0(n32660), .C0(n31034), 
        .Y(n31036) );
  OAI211XL U34137 ( .A0(n33703), .A1(n31037), .B0(n33550), .C0(n31036), .Y(
        n15861) );
  INVXL U34138 ( .A(conv_3[226]), .Y(n31041) );
  OAI211XL U34139 ( .A0(n31039), .A1(conv_3[226]), .B0(n34028), .C0(n31038), 
        .Y(n31040) );
  OAI211XL U34140 ( .A0(n35676), .A1(n31041), .B0(n33550), .C0(n31040), .Y(
        n15872) );
  INVXL U34141 ( .A(conv_3[421]), .Y(n31045) );
  OAI211XL U34142 ( .A0(n31043), .A1(conv_3[421]), .B0(n32181), .C0(n31042), 
        .Y(n31044) );
  OAI211XL U34143 ( .A0(n35778), .A1(n31045), .B0(n33550), .C0(n31044), .Y(
        n15859) );
  INVXL U34144 ( .A(conv_2[211]), .Y(n31051) );
  NAND2XL U34145 ( .A(n31047), .B(n31046), .Y(n31049) );
  NAND2XL U34146 ( .A(n31051), .B(n31049), .Y(n31048) );
  OAI211XL U34147 ( .A0(n31051), .A1(n31049), .B0(n32656), .C0(n31048), .Y(
        n31050) );
  OAI211XL U34148 ( .A0(n35934), .A1(n31051), .B0(n31050), .C0(n35847), .Y(
        n15333) );
  INVXL U34149 ( .A(conv_1[406]), .Y(n31055) );
  OAI211XL U34150 ( .A0(n31053), .A1(conv_1[406]), .B0(n33157), .C0(n31052), 
        .Y(n31054) );
  OAI211XL U34151 ( .A0(n35487), .A1(n31055), .B0(n33067), .C0(n31054), .Y(
        n16057) );
  INVXL U34152 ( .A(conv_2[181]), .Y(n31059) );
  NAND2XL U34153 ( .A(conv_2[181]), .B(n31057), .Y(n31056) );
  OAI211XL U34154 ( .A0(conv_2[181]), .A1(n31057), .B0(n24378), .C0(n31056), 
        .Y(n31058) );
  OAI211XL U34155 ( .A0(n35917), .A1(n31059), .B0(n31058), .C0(n35847), .Y(
        n15335) );
  INVXL U34156 ( .A(conv_3[236]), .Y(n33315) );
  OAI2BB1XL U34157 ( .A0N(conv_3[235]), .A1N(n31061), .B0(n33878), .Y(n33877)
         );
  NAND2XL U34158 ( .A(n33314), .B(n33877), .Y(n31063) );
  AOI211XL U34159 ( .A0(n33315), .A1(n31063), .B0(n34389), .C0(n31062), .Y(
        n31064) );
  AOI2BB1XL U34160 ( .A0N(n33315), .A1N(n35676), .B0(n31064), .Y(n31065) );
  NAND2XL U34161 ( .A(n31065), .B(n35588), .Y(n15587) );
  INVXL U34162 ( .A(conv_2[47]), .Y(n31069) );
  NAND2XL U34163 ( .A(conv_2[47]), .B(n31067), .Y(n31066) );
  OAI211XL U34164 ( .A0(conv_2[47]), .A1(n31067), .B0(n33778), .C0(n31066), 
        .Y(n31068) );
  OAI211XL U34165 ( .A0(n34505), .A1(n31069), .B0(n31068), .C0(n34621), .Y(
        n15308) );
  INVXL U34166 ( .A(weight_1[56]), .Y(n31070) );
  INVXL U34167 ( .A(weight_1[62]), .Y(n31072) );
  OAI22XL U34168 ( .A0(n31084), .A1(n31070), .B0(n31072), .B1(n16647), .Y(
        n14358) );
  INVXL U34169 ( .A(weight_1[50]), .Y(n31074) );
  OAI22XL U34170 ( .A0(n31084), .A1(n31074), .B0(n31070), .B1(n16647), .Y(
        n14357) );
  INVXL U34171 ( .A(weight_1[147]), .Y(n32426) );
  INVXL U34172 ( .A(weight_1[153]), .Y(n32709) );
  OAI22XL U34173 ( .A0(n31084), .A1(n32426), .B0(n32709), .B1(n32840), .Y(
        n14292) );
  INVXL U34174 ( .A(weight_1[213]), .Y(n32440) );
  INVXL U34175 ( .A(weight_1[219]), .Y(n32700) );
  OAI22XL U34176 ( .A0(n31084), .A1(n32440), .B0(n32700), .B1(n32777), .Y(
        n14303) );
  INVXL U34177 ( .A(weight_1[75]), .Y(n31073) );
  INVXL U34178 ( .A(weight_1[81]), .Y(n32425) );
  OAI22XL U34179 ( .A0(n31084), .A1(n31073), .B0(n32425), .B1(n32840), .Y(
        n14280) );
  INVXL U34180 ( .A(weight_1[68]), .Y(n31075) );
  OAI22XL U34181 ( .A0(n31084), .A1(n31072), .B0(n31075), .B1(n16647), .Y(
        n14359) );
  INVXL U34182 ( .A(weight_1[69]), .Y(n32432) );
  OAI22XL U34183 ( .A0(n31084), .A1(n32432), .B0(n31073), .B1(n32840), .Y(
        n14279) );
  INVXL U34184 ( .A(weight_1[44]), .Y(n31076) );
  OAI22XL U34185 ( .A0(n31084), .A1(n31076), .B0(n31074), .B1(n16647), .Y(
        n14356) );
  INVXL U34186 ( .A(weight_1[129]), .Y(n32412) );
  INVXL U34187 ( .A(weight_1[135]), .Y(n32447) );
  OAI22XL U34188 ( .A0(n31084), .A1(n32412), .B0(n32447), .B1(n32840), .Y(
        n14289) );
  INVXL U34189 ( .A(weight_1[74]), .Y(n31079) );
  OAI22XL U34190 ( .A0(n31084), .A1(n31075), .B0(n31079), .B1(n16647), .Y(
        n14360) );
  INVXL U34191 ( .A(weight_1[134]), .Y(n32367) );
  INVXL U34192 ( .A(weight_1[140]), .Y(n32368) );
  OAI22XL U34193 ( .A0(n31084), .A1(n32367), .B0(n32368), .B1(n16647), .Y(
        n14371) );
  INVXL U34194 ( .A(weight_1[38]), .Y(n31078) );
  OAI22XL U34195 ( .A0(n31084), .A1(n31078), .B0(n31076), .B1(n16647), .Y(
        n14355) );
  INVXL U34196 ( .A(weight_1[20]), .Y(n32365) );
  INVXL U34197 ( .A(weight_1[26]), .Y(n31083) );
  OAI22XL U34198 ( .A0(n31084), .A1(n32365), .B0(n31083), .B1(n16647), .Y(
        n14352) );
  INVXL U34199 ( .A(weight_1[86]), .Y(n31080) );
  INVXL U34200 ( .A(weight_1[92]), .Y(n32370) );
  OAI22XL U34201 ( .A0(n31084), .A1(n31080), .B0(n32370), .B1(n16647), .Y(
        n14363) );
  OAI22XL U34202 ( .A0(n31084), .A1(n32387), .B0(n36148), .B1(n16646), .Y(
        n14267) );
  INVXL U34203 ( .A(weight_1[21]), .Y(n32402) );
  INVXL U34204 ( .A(weight_1[27]), .Y(n32766) );
  OAI22XL U34205 ( .A0(n31084), .A1(n32402), .B0(n32766), .B1(n16646), .Y(
        n14271) );
  OAI22XL U34206 ( .A0(n31084), .A1(n32384), .B0(n32385), .B1(n16646), .Y(
        n14260) );
  INVXL U34207 ( .A(weight_1[32]), .Y(n31082) );
  OAI22XL U34208 ( .A0(n31084), .A1(n31082), .B0(n31078), .B1(n16647), .Y(
        n14354) );
  INVXL U34209 ( .A(weight_1[80]), .Y(n31081) );
  OAI22XL U34210 ( .A0(n31084), .A1(n31079), .B0(n31081), .B1(n16647), .Y(
        n14361) );
  OAI22XL U34211 ( .A0(n31084), .A1(n31081), .B0(n31080), .B1(n16647), .Y(
        n14362) );
  OAI22XL U34212 ( .A0(n31084), .A1(n31083), .B0(n31082), .B1(n16647), .Y(
        n14353) );
  INVXL U34213 ( .A(weight_1[98]), .Y(n32369) );
  INVXL U34214 ( .A(weight_1[104]), .Y(n32394) );
  OAI22XL U34215 ( .A0(n31084), .A1(n32369), .B0(n32394), .B1(n16647), .Y(
        n14365) );
  INVXL U34216 ( .A(conv_3[287]), .Y(n31089) );
  ADDFXL U34217 ( .A(conv_3[287]), .B(n31086), .CI(n31085), .CO(n23065), .S(
        n31087) );
  NAND2XL U34218 ( .A(n32611), .B(n31087), .Y(n31088) );
  OAI211XL U34219 ( .A0(n35726), .A1(n31089), .B0(n31088), .C0(n35566), .Y(
        n15832) );
  INVXL U34220 ( .A(conv_2[166]), .Y(n31093) );
  OAI211XL U34221 ( .A0(n31091), .A1(conv_2[166]), .B0(n33157), .C0(n31090), 
        .Y(n31092) );
  OAI211XL U34222 ( .A0(n34589), .A1(n31093), .B0(n35847), .C0(n31092), .Y(
        n15336) );
  INVXL U34223 ( .A(conv_2[196]), .Y(n31097) );
  OAI211XL U34224 ( .A0(n31095), .A1(conv_2[196]), .B0(n32611), .C0(n31094), 
        .Y(n31096) );
  OAI211XL U34225 ( .A0(n35931), .A1(n31097), .B0(n35847), .C0(n31096), .Y(
        n15334) );
  INVXL U34226 ( .A(conv_2[226]), .Y(n31101) );
  OAI211XL U34227 ( .A0(n31099), .A1(conv_2[226]), .B0(n34028), .C0(n31098), 
        .Y(n31100) );
  OAI211XL U34228 ( .A0(n34458), .A1(n31101), .B0(n35847), .C0(n31100), .Y(
        n15332) );
  INVXL U34229 ( .A(conv_2[32]), .Y(n31107) );
  NOR2BXL U34230 ( .AN(n31103), .B(n31102), .Y(n31105) );
  NAND2XL U34231 ( .A(conv_2[32]), .B(n31105), .Y(n31104) );
  OAI211XL U34232 ( .A0(conv_2[32]), .A1(n31105), .B0(n33778), .C0(n31104), 
        .Y(n31106) );
  OAI211XL U34233 ( .A0(n35865), .A1(n31107), .B0(n34621), .C0(n31106), .Y(
        n15309) );
  OAI2BB1XL U34234 ( .A0N(n36020), .A1N(n31108), .B0(n35826), .Y(n31109) );
  AOI32XL U34235 ( .A0(n34742), .A1(n31109), .A2(n33530), .B0(conv_3[480]), 
        .B1(n31109), .Y(n31110) );
  NAND2XL U34236 ( .A(n34755), .B(n31110), .Y(n15891) );
  OAI2BB1XL U34237 ( .A0N(conv_1[205]), .A1N(n35378), .B0(n34060), .Y(n35386)
         );
  NAND4XL U34238 ( .A(conv_1[206]), .B(conv_1[207]), .C(n34060), .D(n35386), 
        .Y(n33118) );
  OAI21XL U34239 ( .A0(conv_1[205]), .A1(n35377), .B0(n35379), .Y(n35385) );
  INVXL U34240 ( .A(conv_1[207]), .Y(n34064) );
  NAND3XL U34241 ( .A(n35387), .B(n35379), .C(n34064), .Y(n33117) );
  NAND2XL U34242 ( .A(n33118), .B(n33117), .Y(n31115) );
  NAND2XL U34243 ( .A(conv_1[208]), .B(n31115), .Y(n31114) );
  OAI211XL U34244 ( .A0(conv_1[208]), .A1(n31115), .B0(n33712), .C0(n31114), 
        .Y(n31116) );
  OAI211XL U34245 ( .A0(n35384), .A1(n33116), .B0(n16652), .C0(n31116), .Y(
        n16255) );
  NAND2XL U34246 ( .A(n33097), .B(n33096), .Y(n33095) );
  OAI21XL U34247 ( .A0(n33097), .A1(n33096), .B0(n33095), .Y(n31119) );
  NAND2XL U34248 ( .A(conv_2[238]), .B(n31119), .Y(n31118) );
  OAI211XL U34249 ( .A0(conv_2[238]), .A1(n31119), .B0(n34028), .C0(n31118), 
        .Y(n31120) );
  OAI211XL U34250 ( .A0(n34458), .A1(n33094), .B0(n35859), .C0(n31120), .Y(
        n15045) );
  NAND4XL U34251 ( .A(conv_2[221]), .B(conv_2[222]), .C(n31121), .D(n35936), 
        .Y(n33264) );
  NAND3XL U34252 ( .A(n35937), .B(n33770), .C(n31122), .Y(n33263) );
  AOI22XL U34253 ( .A0(conv_2[223]), .A1(n33264), .B0(n33263), .B1(n33267), 
        .Y(n31124) );
  NAND2XL U34254 ( .A(conv_2[224]), .B(n31124), .Y(n31123) );
  OAI211XL U34255 ( .A0(conv_2[224]), .A1(n31124), .B0(n33982), .C0(n31123), 
        .Y(n31125) );
  OAI211XL U34256 ( .A0(n33853), .A1(n31126), .B0(n35859), .C0(n31125), .Y(
        n15054) );
  OAI21XL U34257 ( .A0(conv_1[235]), .A1(n31127), .B0(n35404), .Y(n31129) );
  AND2X1 U34258 ( .A(n31130), .B(n31129), .Y(n34274) );
  AOI31XL U34259 ( .A0(n36020), .A1(n34274), .A2(n34275), .B0(n35549), .Y(
        n31132) );
  OAI2BB1XL U34260 ( .A0N(n31129), .A1N(n34275), .B0(n34028), .Y(n31131) );
  AOI32XL U34261 ( .A0(n35408), .A1(n31132), .A2(n31131), .B0(n31130), .B1(
        n31132), .Y(n16227) );
  INVXL U34262 ( .A(conv_2[58]), .Y(n33102) );
  NAND4XL U34263 ( .A(conv_2[56]), .B(conv_2[57]), .C(n31134), .D(n31133), .Y(
        n33104) );
  NAND3XL U34264 ( .A(n31137), .B(n31136), .C(n31135), .Y(n33103) );
  NAND2XL U34265 ( .A(n33104), .B(n33103), .Y(n31139) );
  NAND2XL U34266 ( .A(conv_2[58]), .B(n31139), .Y(n31138) );
  OAI211XL U34267 ( .A0(conv_2[58]), .A1(n31139), .B0(n16657), .C0(n31138), 
        .Y(n31140) );
  OAI211XL U34268 ( .A0(n34505), .A1(n33102), .B0(n33815), .C0(n31140), .Y(
        n15165) );
  INVXL U34269 ( .A(conv_3[535]), .Y(n31146) );
  AOI2BB1XL U34270 ( .A0N(n33719), .A1N(n31142), .B0(n31141), .Y(n31144) );
  NAND2XL U34271 ( .A(conv_3[535]), .B(n31144), .Y(n31143) );
  OAI211XL U34272 ( .A0(conv_3[535]), .A1(n31144), .B0(n24499), .C0(n31143), 
        .Y(n31145) );
  OAI211XL U34273 ( .A0(n31191), .A1(n31146), .B0(n16649), .C0(n31145), .Y(
        n15388) );
  NAND2XL U34274 ( .A(conv_3[519]), .B(n31150), .Y(n31149) );
  OAI211XL U34275 ( .A0(conv_3[519]), .A1(n31150), .B0(n34666), .C0(n31149), 
        .Y(n31151) );
  OAI211XL U34276 ( .A0(n33303), .A1(n31152), .B0(n16649), .C0(n31151), .Y(
        n15399) );
  INVXL U34277 ( .A(conv_3[522]), .Y(n31157) );
  NAND2XL U34278 ( .A(n31292), .B(conv_3[521]), .Y(n31153) );
  OAI32XL U34279 ( .A0(n31291), .A1(n31292), .A2(conv_3[521]), .B0(n31180), 
        .B1(n31153), .Y(n31155) );
  NAND2XL U34280 ( .A(conv_3[522]), .B(n31155), .Y(n31154) );
  OAI211XL U34281 ( .A0(conv_3[522]), .A1(n31155), .B0(n16657), .C0(n31154), 
        .Y(n31156) );
  OAI211XL U34282 ( .A0(n33303), .A1(n31157), .B0(n16649), .C0(n31156), .Y(
        n15396) );
  INVXL U34283 ( .A(conv_3[9]), .Y(n31161) );
  NAND2XL U34284 ( .A(conv_3[9]), .B(n31159), .Y(n31158) );
  OAI211XL U34285 ( .A0(conv_3[9]), .A1(n31159), .B0(n33157), .C0(n31158), .Y(
        n31160) );
  OAI211XL U34286 ( .A0(n34383), .A1(n31161), .B0(n33468), .C0(n31160), .Y(
        n15739) );
  OAI32XL U34287 ( .A0(n31291), .A1(n31173), .A2(conv_3[516]), .B0(n31180), 
        .B1(n31162), .Y(n31164) );
  NAND2XL U34288 ( .A(conv_3[517]), .B(n31164), .Y(n31163) );
  OAI211XL U34289 ( .A0(conv_3[517]), .A1(n31164), .B0(n24499), .C0(n31163), 
        .Y(n31165) );
  OAI211XL U34290 ( .A0(n33303), .A1(n31166), .B0(n16649), .C0(n31165), .Y(
        n15401) );
  AOI32XL U34291 ( .A0(conv_3[536]), .A1(n31167), .A2(n31185), .B0(n33719), 
        .B1(n31167), .Y(n31169) );
  NAND2XL U34292 ( .A(n31171), .B(n31169), .Y(n31168) );
  OAI211XL U34293 ( .A0(n31171), .A1(n31169), .B0(n34666), .C0(n31168), .Y(
        n31170) );
  OAI211XL U34294 ( .A0(n31191), .A1(n31171), .B0(n16649), .C0(n31170), .Y(
        n15386) );
  AOI21XL U34295 ( .A0(n31173), .A1(n31180), .B0(n31172), .Y(n31175) );
  NAND2XL U34296 ( .A(conv_3[516]), .B(n31175), .Y(n31174) );
  OAI211XL U34297 ( .A0(conv_3[516]), .A1(n31175), .B0(n32611), .C0(n31174), 
        .Y(n31176) );
  OAI211XL U34298 ( .A0(n33303), .A1(n31177), .B0(n33468), .C0(n31176), .Y(
        n15402) );
  OAI21XL U34299 ( .A0(n31180), .A1(n31179), .B0(n31178), .Y(n31182) );
  NAND2XL U34300 ( .A(n31184), .B(n31182), .Y(n31181) );
  OAI211XL U34301 ( .A0(n31184), .A1(n31182), .B0(n31735), .C0(n31181), .Y(
        n31183) );
  OAI211XL U34302 ( .A0(n33303), .A1(n31184), .B0(n16649), .C0(n31183), .Y(
        n15400) );
  NAND2XL U34303 ( .A(n31186), .B(n31185), .Y(n31188) );
  NAND2XL U34304 ( .A(n31190), .B(n31188), .Y(n31187) );
  OAI211XL U34305 ( .A0(n31190), .A1(n31188), .B0(n32656), .C0(n31187), .Y(
        n31189) );
  OAI211XL U34306 ( .A0(n31191), .A1(n31190), .B0(n33468), .C0(n31189), .Y(
        n15387) );
  AOI22XL U34307 ( .A0(conv_3[8]), .A1(n34379), .B0(n32996), .B1(n31196), .Y(
        n31193) );
  NAND2XL U34308 ( .A(n31194), .B(n31193), .Y(n31192) );
  OAI211XL U34309 ( .A0(n31194), .A1(n31193), .B0(n33157), .C0(n31192), .Y(
        n31195) );
  OAI211XL U34310 ( .A0(n34383), .A1(n31196), .B0(n16649), .C0(n31195), .Y(
        n15740) );
  NAND2XL U34311 ( .A(n31198), .B(n31197), .Y(n31216) );
  OAI2BB1XL U34312 ( .A0N(conv_3[54]), .A1N(n31199), .B0(n32178), .Y(n31217)
         );
  OAI2BB1XL U34313 ( .A0N(n33824), .A1N(n31216), .B0(n31217), .Y(n31201) );
  NAND2XL U34314 ( .A(n31203), .B(n31201), .Y(n31200) );
  OAI211XL U34315 ( .A0(n31203), .A1(n31201), .B0(n33982), .C0(n31200), .Y(
        n31202) );
  OAI211XL U34316 ( .A0(n34392), .A1(n31203), .B0(n16649), .C0(n31202), .Y(
        n15708) );
  INVXL U34317 ( .A(conv_3[52]), .Y(n31209) );
  AOI2BB1XL U34318 ( .A0N(n33824), .A1N(n31205), .B0(n31204), .Y(n31207) );
  NAND2XL U34319 ( .A(conv_3[52]), .B(n31207), .Y(n31206) );
  OAI211XL U34320 ( .A0(conv_3[52]), .A1(n31207), .B0(n35336), .C0(n31206), 
        .Y(n31208) );
  OAI211XL U34321 ( .A0(n34392), .A1(n31209), .B0(n16649), .C0(n31208), .Y(
        n15711) );
  AOI21XL U34322 ( .A0(n33824), .A1(n31211), .B0(n31210), .Y(n31213) );
  NAND2XL U34323 ( .A(conv_3[51]), .B(n31213), .Y(n31212) );
  OAI211XL U34324 ( .A0(conv_3[51]), .A1(n31213), .B0(n16657), .C0(n31212), 
        .Y(n31214) );
  OAI211XL U34325 ( .A0(n34392), .A1(n31215), .B0(n33468), .C0(n31214), .Y(
        n15712) );
  INVXL U34326 ( .A(conv_3[56]), .Y(n31221) );
  AOI21XL U34327 ( .A0(conv_3[55]), .A1(n31217), .B0(n33824), .Y(n32177) );
  NAND2XL U34328 ( .A(conv_3[56]), .B(n31219), .Y(n31218) );
  OAI211XL U34329 ( .A0(conv_3[56]), .A1(n31219), .B0(n16656), .C0(n31218), 
        .Y(n31220) );
  OAI211XL U34330 ( .A0(n34392), .A1(n31221), .B0(n33468), .C0(n31220), .Y(
        n15707) );
  NAND3XL U34331 ( .A(conv_3[42]), .B(n31239), .C(n35591), .Y(n31299) );
  OR3XL U34332 ( .A(n31239), .B(conv_3[42]), .C(n35591), .Y(n31298) );
  NAND2XL U34333 ( .A(n31299), .B(n31298), .Y(n31224) );
  NAND2XL U34334 ( .A(conv_3[43]), .B(n31224), .Y(n31223) );
  OAI211XL U34335 ( .A0(conv_3[43]), .A1(n31224), .B0(n30090), .C0(n31223), 
        .Y(n31225) );
  OAI211XL U34336 ( .A0(n35594), .A1(n31297), .B0(n16649), .C0(n31225), .Y(
        n15715) );
  AOI2BB1XL U34337 ( .A0N(n33449), .A1N(n31227), .B0(n31226), .Y(n31229) );
  NAND2XL U34338 ( .A(conv_3[39]), .B(n31229), .Y(n31228) );
  OAI211XL U34339 ( .A0(conv_3[39]), .A1(n31229), .B0(n36020), .C0(n31228), 
        .Y(n31230) );
  OAI211XL U34340 ( .A0(n35594), .A1(n31231), .B0(n33468), .C0(n31230), .Y(
        n15719) );
  NAND2XL U34341 ( .A(conv_3[40]), .B(n31235), .Y(n31234) );
  OAI211XL U34342 ( .A0(conv_3[40]), .A1(n31235), .B0(n27932), .C0(n31234), 
        .Y(n31236) );
  OAI211XL U34343 ( .A0(n35594), .A1(n31237), .B0(n16649), .C0(n31236), .Y(
        n15718) );
  INVXL U34344 ( .A(conv_3[42]), .Y(n31243) );
  AOI21XL U34345 ( .A0(n31239), .A1(n33449), .B0(n31238), .Y(n31241) );
  NAND2XL U34346 ( .A(conv_3[42]), .B(n31241), .Y(n31240) );
  OAI211XL U34347 ( .A0(conv_3[42]), .A1(n31241), .B0(n30090), .C0(n31240), 
        .Y(n31242) );
  OAI211XL U34348 ( .A0(n35594), .A1(n31243), .B0(n16649), .C0(n31242), .Y(
        n15716) );
  AOI21XL U34349 ( .A0(n35591), .A1(n31245), .B0(n31244), .Y(n31247) );
  NAND2XL U34350 ( .A(conv_3[36]), .B(n31247), .Y(n31246) );
  OAI211XL U34351 ( .A0(conv_3[36]), .A1(n31247), .B0(n33157), .C0(n31246), 
        .Y(n31248) );
  OAI211XL U34352 ( .A0(n35594), .A1(n31249), .B0(n33468), .C0(n31248), .Y(
        n15722) );
  AOI2BB1XL U34353 ( .A0N(n33002), .A1N(n31257), .B0(n31258), .Y(n31254) );
  NAND2XL U34354 ( .A(conv_3[25]), .B(n31254), .Y(n31253) );
  OAI211XL U34355 ( .A0(conv_3[25]), .A1(n31254), .B0(n33157), .C0(n31253), 
        .Y(n31255) );
  OAI211XL U34356 ( .A0(n35576), .A1(n31256), .B0(n33468), .C0(n31255), .Y(
        n15728) );
  INVXL U34357 ( .A(conv_3[27]), .Y(n31305) );
  OAI2BB1XL U34358 ( .A0N(conv_3[25]), .A1N(n31257), .B0(n31304), .Y(n35578)
         );
  OAI21XL U34359 ( .A0(conv_3[25]), .A1(n31258), .B0(n33002), .Y(n35577) );
  AOI32XL U34360 ( .A0(conv_3[26]), .A1(n31304), .A2(n35578), .B0(n33002), 
        .B1(n35579), .Y(n31260) );
  NAND2XL U34361 ( .A(n31305), .B(n31260), .Y(n31259) );
  OAI211XL U34362 ( .A0(n31305), .A1(n31260), .B0(n33157), .C0(n31259), .Y(
        n31261) );
  OAI211XL U34363 ( .A0(n35576), .A1(n31305), .B0(n16649), .C0(n31261), .Y(
        n15726) );
  AOI221XL U34364 ( .A0(conv_3[21]), .A1(n33002), .B0(n31274), .B1(n33002), 
        .C0(n31262), .Y(n31264) );
  NAND2XL U34365 ( .A(conv_3[22]), .B(n31264), .Y(n31263) );
  OAI211XL U34366 ( .A0(conv_3[22]), .A1(n31264), .B0(n33157), .C0(n31263), 
        .Y(n31265) );
  OAI211XL U34367 ( .A0(n35576), .A1(n31266), .B0(n16649), .C0(n31265), .Y(
        n15731) );
  OAI21XL U34368 ( .A0(n33002), .A1(n31268), .B0(n31267), .Y(n31270) );
  NAND2XL U34369 ( .A(n31272), .B(n31270), .Y(n31269) );
  OAI211XL U34370 ( .A0(n31272), .A1(n31270), .B0(n33157), .C0(n31269), .Y(
        n31271) );
  OAI211XL U34371 ( .A0(n35576), .A1(n31272), .B0(n33468), .C0(n31271), .Y(
        n15730) );
  AOI21XL U34372 ( .A0(n31274), .A1(n33002), .B0(n31273), .Y(n31276) );
  NAND2XL U34373 ( .A(conv_3[21]), .B(n31276), .Y(n31275) );
  OAI211XL U34374 ( .A0(conv_3[21]), .A1(n31276), .B0(n33157), .C0(n31275), 
        .Y(n31277) );
  OAI211XL U34375 ( .A0(n35576), .A1(n31278), .B0(n33468), .C0(n31277), .Y(
        n15732) );
  INVXL U34376 ( .A(conv_1[399]), .Y(n35473) );
  NAND2XL U34377 ( .A(conv_1[398]), .B(n31279), .Y(n35470) );
  OAI2BB1XL U34378 ( .A0N(conv_1[400]), .A1N(n33653), .B0(n35471), .Y(n35479)
         );
  AOI32XL U34379 ( .A0(conv_1[401]), .A1(n35471), .A2(n35479), .B0(n33654), 
        .B1(n35480), .Y(n31282) );
  NAND2XL U34380 ( .A(n33269), .B(n31282), .Y(n31281) );
  OAI211XL U34381 ( .A0(n33269), .A1(n31282), .B0(n32052), .C0(n31281), .Y(
        n31283) );
  OAI211XL U34382 ( .A0(n35477), .A1(n33269), .B0(n34544), .C0(n31283), .Y(
        n16061) );
  AOI22XL U34383 ( .A0(conv_3[538]), .A1(n31286), .B0(n31285), .B1(n31284), 
        .Y(n31288) );
  NAND2XL U34384 ( .A(conv_3[539]), .B(n31288), .Y(n31287) );
  OAI211XL U34385 ( .A0(conv_3[539]), .A1(n31288), .B0(n33778), .C0(n31287), 
        .Y(n31289) );
  OAI211XL U34386 ( .A0(n33853), .A1(n31290), .B0(n33468), .C0(n31289), .Y(
        n15384) );
  NAND4XL U34387 ( .A(conv_3[522]), .B(conv_3[521]), .C(n31292), .D(n31291), 
        .Y(n33302) );
  INVXL U34388 ( .A(conv_3[523]), .Y(n33306) );
  AOI22XL U34389 ( .A0(conv_3[523]), .A1(n33302), .B0(n33301), .B1(n33306), 
        .Y(n31294) );
  NAND2XL U34390 ( .A(conv_3[524]), .B(n31294), .Y(n31293) );
  OAI211XL U34391 ( .A0(conv_3[524]), .A1(n31294), .B0(n34666), .C0(n31293), 
        .Y(n31295) );
  OAI211XL U34392 ( .A0(n34520), .A1(n31296), .B0(n33468), .C0(n31295), .Y(
        n15394) );
  AOI22XL U34393 ( .A0(conv_3[43]), .A1(n31299), .B0(n31298), .B1(n31297), .Y(
        n31301) );
  NAND2XL U34394 ( .A(conv_3[44]), .B(n31301), .Y(n31300) );
  OAI211XL U34395 ( .A0(conv_3[44]), .A1(n31301), .B0(n35336), .C0(n31300), 
        .Y(n31302) );
  OAI211XL U34396 ( .A0(n34789), .A1(n31303), .B0(n16649), .C0(n31302), .Y(
        n15714) );
  NAND4XL U34397 ( .A(conv_3[26]), .B(conv_3[27]), .C(n31304), .D(n35578), .Y(
        n34411) );
  NAND3XL U34398 ( .A(n35579), .B(n33002), .C(n31305), .Y(n34410) );
  AOI22XL U34399 ( .A0(conv_3[28]), .A1(n34411), .B0(n34410), .B1(n34414), .Y(
        n31307) );
  NAND2XL U34400 ( .A(conv_3[29]), .B(n31307), .Y(n31306) );
  OAI211XL U34401 ( .A0(conv_3[29]), .A1(n31307), .B0(n33157), .C0(n31306), 
        .Y(n31308) );
  OAI211XL U34402 ( .A0(n34789), .A1(n31309), .B0(n33468), .C0(n31308), .Y(
        n15724) );
  INVXL U34403 ( .A(conv_2[208]), .Y(n33034) );
  NAND3XL U34404 ( .A(conv_2[207]), .B(n31310), .C(n35928), .Y(n33036) );
  OR3XL U34405 ( .A(n31310), .B(conv_2[207]), .C(n35928), .Y(n33035) );
  NAND2XL U34406 ( .A(n33036), .B(n33035), .Y(n31312) );
  OAI21XL U34407 ( .A0(n36009), .A1(n31312), .B0(n35931), .Y(n31311) );
  AOI32XL U34408 ( .A0(n36020), .A1(n33034), .A2(n31312), .B0(conv_2[208]), 
        .B1(n31311), .Y(n31313) );
  NAND2XL U34409 ( .A(n31313), .B(n35859), .Y(n15065) );
  INVXL U34410 ( .A(weight_1[31]), .Y(n32350) );
  INVXL U34411 ( .A(weight_1[37]), .Y(n31314) );
  OAI22XL U34412 ( .A0(n31084), .A1(n32350), .B0(n31314), .B1(n26910), .Y(
        n14435) );
  INVXL U34413 ( .A(weight_1[103]), .Y(n32356) );
  INVXL U34414 ( .A(weight_1[109]), .Y(n32354) );
  OAI22XL U34415 ( .A0(n31071), .A1(n32356), .B0(n32354), .B1(n26910), .Y(
        n14447) );
  INVXL U34416 ( .A(weight_1[67]), .Y(n32683) );
  INVXL U34417 ( .A(weight_1[73]), .Y(n32686) );
  OAI22XL U34418 ( .A0(n32491), .A1(n32683), .B0(n32686), .B1(n26910), .Y(
        n14441) );
  INVXL U34419 ( .A(weight_1[43]), .Y(n32681) );
  OAI22XL U34420 ( .A0(n16650), .A1(n31314), .B0(n32681), .B1(n26910), .Y(
        n14436) );
  OAI22XL U34421 ( .A0(n16650), .A1(n32355), .B0(n32679), .B1(n26910), .Y(
        n14427) );
  INVXL U34422 ( .A(weight_1[60]), .Y(n31316) );
  INVXL U34423 ( .A(weight_1[66]), .Y(n31327) );
  OAI22XL U34424 ( .A0(n31071), .A1(n31316), .B0(n31327), .B1(n32840), .Y(
        n14521) );
  INVXL U34425 ( .A(weight_1[422]), .Y(n32366) );
  OAI22XL U34426 ( .A0(n32491), .A1(n32366), .B0(n32390), .B1(n16646), .Y(
        n14419) );
  INVXL U34427 ( .A(weight_1[48]), .Y(n32737) );
  INVXL U34428 ( .A(weight_1[54]), .Y(n31317) );
  OAI22XL U34429 ( .A0(n16645), .A1(n32737), .B0(n31317), .B1(n16648), .Y(
        n14519) );
  INVXL U34430 ( .A(weight_1[409]), .Y(n32696) );
  INVXL U34431 ( .A(weight_1[415]), .Y(n32423) );
  OAI22XL U34432 ( .A0(n16650), .A1(n32696), .B0(n32423), .B1(n16648), .Y(
        n14498) );
  INVXL U34433 ( .A(weight_1[84]), .Y(n31320) );
  INVXL U34434 ( .A(weight_1[90]), .Y(n31315) );
  OAI22XL U34435 ( .A0(n32491), .A1(n31320), .B0(n31315), .B1(n16646), .Y(
        n14525) );
  INVXL U34436 ( .A(weight_1[96]), .Y(n31323) );
  OAI22XL U34437 ( .A0(n16645), .A1(n31315), .B0(n31323), .B1(n16647), .Y(
        n14526) );
  OAI22XL U34438 ( .A0(n31071), .A1(n31317), .B0(n31316), .B1(n26910), .Y(
        n14520) );
  INVXL U34439 ( .A(weight_1[72]), .Y(n31326) );
  INVXL U34440 ( .A(weight_1[78]), .Y(n31321) );
  OAI22XL U34441 ( .A0(n32491), .A1(n31326), .B0(n31321), .B1(n26910), .Y(
        n14523) );
  INVXL U34442 ( .A(weight_1[12]), .Y(n32723) );
  INVXL U34443 ( .A(weight_1[18]), .Y(n32411) );
  OAI22XL U34444 ( .A0(n16650), .A1(n32723), .B0(n32411), .B1(n26910), .Y(
        n14513) );
  INVXL U34445 ( .A(weight_1[120]), .Y(n31319) );
  OAI22XL U34446 ( .A0(n16645), .A1(n31319), .B0(n31318), .B1(n16648), .Y(
        n14531) );
  INVXL U34447 ( .A(weight_1[114]), .Y(n31324) );
  OAI22XL U34448 ( .A0(n32491), .A1(n31324), .B0(n31319), .B1(n32840), .Y(
        n14530) );
  OAI22XL U34449 ( .A0(n16650), .A1(n31321), .B0(n31320), .B1(n16646), .Y(
        n14524) );
  INVXL U34450 ( .A(weight_1[102]), .Y(n31322) );
  INVXL U34451 ( .A(weight_1[108]), .Y(n31325) );
  OAI22XL U34452 ( .A0(n16650), .A1(n31322), .B0(n31325), .B1(n26910), .Y(
        n14528) );
  OAI22XL U34453 ( .A0(n26906), .A1(n31323), .B0(n31322), .B1(n16647), .Y(
        n14527) );
  OAI22XL U34454 ( .A0(n16650), .A1(n31325), .B0(n31324), .B1(n26910), .Y(
        n14529) );
  OAI22XL U34455 ( .A0(n31077), .A1(n31327), .B0(n31326), .B1(n32777), .Y(
        n14522) );
  OAI22XL U34456 ( .A0(n31084), .A1(n31328), .B0(n32419), .B1(n16648), .Y(
        n14505) );
  OAI22XL U34457 ( .A0(n32491), .A1(n32727), .B0(n31328), .B1(n16648), .Y(
        n14504) );
  INVXL U34458 ( .A(conv_3[360]), .Y(n31332) );
  OAI211XL U34459 ( .A0(conv_3[360]), .A1(n31330), .B0(n33912), .C0(n31329), 
        .Y(n31331) );
  OAI211XL U34460 ( .A0(n35764), .A1(n31332), .B0(n31331), .C0(n34755), .Y(
        n15899) );
  NAND4XL U34461 ( .A(conv_1[101]), .B(conv_1[102]), .C(n31334), .D(n31333), 
        .Y(n31356) );
  NAND3XL U34462 ( .A(n31337), .B(n31336), .C(n31335), .Y(n31355) );
  INVXL U34463 ( .A(conv_1[103]), .Y(n31360) );
  AOI22XL U34464 ( .A0(conv_1[103]), .A1(n31356), .B0(n31355), .B1(n31360), 
        .Y(n31339) );
  NAND2XL U34465 ( .A(conv_1[104]), .B(n31339), .Y(n31338) );
  OAI211XL U34466 ( .A0(conv_1[104]), .A1(n31339), .B0(n34028), .C0(n31338), 
        .Y(n31340) );
  OAI32XL U34467 ( .A0(n31344), .A1(conv_1[113]), .A2(n31343), .B0(n34557), 
        .B1(n31342), .Y(n31346) );
  NAND2XL U34468 ( .A(conv_1[114]), .B(n31346), .Y(n31345) );
  OAI211XL U34469 ( .A0(conv_1[114]), .A1(n31346), .B0(n32611), .C0(n31345), 
        .Y(n31347) );
  OAI211XL U34470 ( .A0(n35330), .A1(n31348), .B0(n34682), .C0(n31347), .Y(
        n16349) );
  NAND2XL U34471 ( .A(conv_1[111]), .B(n31352), .Y(n31351) );
  OAI211XL U34472 ( .A0(conv_1[111]), .A1(n31352), .B0(n33778), .C0(n31351), 
        .Y(n31353) );
  OAI211XL U34473 ( .A0(n35330), .A1(n31354), .B0(n16652), .C0(n31353), .Y(
        n16352) );
  NAND2XL U34474 ( .A(n31356), .B(n31355), .Y(n31358) );
  NAND2XL U34475 ( .A(conv_1[103]), .B(n31358), .Y(n31357) );
  OAI211XL U34476 ( .A0(conv_1[103]), .A1(n31358), .B0(n32656), .C0(n31357), 
        .Y(n31359) );
  OAI211XL U34477 ( .A0(n31361), .A1(n31360), .B0(n34689), .C0(n31359), .Y(
        n16360) );
  INVXL U34478 ( .A(conv_1[373]), .Y(n33128) );
  OAI2BB1XL U34479 ( .A0N(conv_1[370]), .A1N(n31362), .B0(n31363), .Y(n34306)
         );
  NAND4XL U34480 ( .A(conv_1[371]), .B(conv_1[372]), .C(n31363), .D(n34306), 
        .Y(n33130) );
  INVXL U34481 ( .A(conv_1[371]), .Y(n34287) );
  OAI21XL U34482 ( .A0(conv_1[370]), .A1(n31364), .B0(n35455), .Y(n34283) );
  NAND2XL U34483 ( .A(n34287), .B(n34283), .Y(n31365) );
  NAND3XL U34484 ( .A(n35455), .B(n34311), .C(n34307), .Y(n33129) );
  NAND2XL U34485 ( .A(n33130), .B(n33129), .Y(n31367) );
  NAND2XL U34486 ( .A(conv_1[373]), .B(n31367), .Y(n31366) );
  OAI211XL U34487 ( .A0(conv_1[373]), .A1(n31367), .B0(n16657), .C0(n31366), 
        .Y(n31368) );
  OAI211XL U34488 ( .A0(n35458), .A1(n33128), .B0(n34544), .C0(n31368), .Y(
        n16090) );
  INVXL U34489 ( .A(conv_1[108]), .Y(n31375) );
  AOI21XL U34490 ( .A0(n31371), .A1(n31370), .B0(n31369), .Y(n31373) );
  NAND2XL U34491 ( .A(conv_1[108]), .B(n31373), .Y(n31372) );
  OAI211XL U34492 ( .A0(conv_1[108]), .A1(n31373), .B0(n33982), .C0(n31372), 
        .Y(n31374) );
  OAI211XL U34493 ( .A0(n35330), .A1(n31375), .B0(n31374), .C0(n32867), .Y(
        n16355) );
  OAI211XL U34494 ( .A0(n31377), .A1(conv_3[465]), .B0(n33912), .C0(n31376), 
        .Y(n31378) );
  OAI211XL U34495 ( .A0(n35813), .A1(n31379), .B0(n34755), .C0(n31378), .Y(
        n15892) );
  INVXL U34496 ( .A(conv_3[495]), .Y(n31383) );
  OAI211XL U34497 ( .A0(n31381), .A1(conv_3[495]), .B0(n33912), .C0(n31380), 
        .Y(n31382) );
  OAI211XL U34498 ( .A0(n35841), .A1(n31383), .B0(n34755), .C0(n31382), .Y(
        n15890) );
  INVXL U34499 ( .A(conv_3[386]), .Y(n31390) );
  NAND2XL U34500 ( .A(n34164), .B(n31502), .Y(n31501) );
  NAND2XL U34501 ( .A(n31506), .B(n31501), .Y(n31461) );
  INVXL U34502 ( .A(n34164), .Y(n32200) );
  AOI31XL U34503 ( .A0(conv_3[385]), .A1(conv_3[384]), .A2(n31502), .B0(n34164), .Y(n32198) );
  NAND2XL U34504 ( .A(conv_3[386]), .B(n31388), .Y(n31387) );
  OAI211XL U34505 ( .A0(conv_3[386]), .A1(n31388), .B0(n30090), .C0(n31387), 
        .Y(n31389) );
  OAI211XL U34506 ( .A0(n34168), .A1(n31390), .B0(n16649), .C0(n31389), .Y(
        n15487) );
  INVXL U34507 ( .A(conv_3[351]), .Y(n31397) );
  INVXL U34508 ( .A(n32130), .Y(n33752) );
  AND2XL U34509 ( .A(n32130), .B(n31393), .Y(n31479) );
  AOI2BB1XL U34510 ( .A0N(n33752), .A1N(n31449), .B0(n31450), .Y(n31395) );
  NAND2XL U34511 ( .A(conv_3[351]), .B(n31395), .Y(n31394) );
  OAI211XL U34512 ( .A0(conv_3[351]), .A1(n31395), .B0(n33157), .C0(n31394), 
        .Y(n31396) );
  OAI211XL U34513 ( .A0(n34746), .A1(n31397), .B0(n16649), .C0(n31396), .Y(
        n15512) );
  NAND2XL U34514 ( .A(conv_3[125]), .B(n31401), .Y(n31400) );
  OAI211XL U34515 ( .A0(conv_3[125]), .A1(n31401), .B0(n16657), .C0(n31400), 
        .Y(n31402) );
  OAI211XL U34516 ( .A0(n35626), .A1(n31403), .B0(n33468), .C0(n31402), .Y(
        n15663) );
  INVXL U34517 ( .A(conv_3[308]), .Y(n31411) );
  INVXL U34518 ( .A(conv_3[307]), .Y(n35735) );
  INVXL U34519 ( .A(n35732), .Y(n33109) );
  AOI2BB1XL U34520 ( .A0N(conv_3[307]), .A1N(n35733), .B0(n33109), .Y(n31407)
         );
  AOI2BB1XL U34521 ( .A0N(n35732), .A1N(n31496), .B0(n31407), .Y(n31409) );
  NAND2XL U34522 ( .A(conv_3[308]), .B(n31409), .Y(n31408) );
  OAI211XL U34523 ( .A0(conv_3[308]), .A1(n31409), .B0(n16656), .C0(n31408), 
        .Y(n31410) );
  OAI211XL U34524 ( .A0(n35736), .A1(n31411), .B0(n33468), .C0(n31410), .Y(
        n15540) );
  INVXL U34525 ( .A(conv_3[128]), .Y(n31417) );
  AOI2BB1XL U34526 ( .A0N(n35622), .A1N(n31413), .B0(n31412), .Y(n31415) );
  NAND2XL U34527 ( .A(conv_3[128]), .B(n31415), .Y(n31414) );
  OAI211XL U34528 ( .A0(conv_3[128]), .A1(n31415), .B0(n24378), .C0(n31414), 
        .Y(n31416) );
  OAI211XL U34529 ( .A0(n35626), .A1(n31417), .B0(n33468), .C0(n31416), .Y(
        n15660) );
  INVXL U34530 ( .A(conv_3[72]), .Y(n31425) );
  OAI31XL U34531 ( .A0(conv_3[67]), .A1(n35600), .A2(conv_3[68]), .B0(n35599), 
        .Y(n31473) );
  INVXL U34532 ( .A(n35599), .Y(n32163) );
  INVXL U34533 ( .A(conv_3[68]), .Y(n31495) );
  NOR2X1 U34534 ( .A(n31491), .B(n31495), .Y(n31474) );
  AOI21X1 U34535 ( .A0(n31474), .A1(conv_3[69]), .B0(n35599), .Y(n31431) );
  AOI21XL U34536 ( .A0(n32164), .A1(n35599), .B0(n31421), .Y(n31423) );
  NAND2XL U34537 ( .A(conv_3[72]), .B(n31423), .Y(n31422) );
  OAI211XL U34538 ( .A0(conv_3[72]), .A1(n31423), .B0(n31735), .C0(n31422), 
        .Y(n31424) );
  OAI211XL U34539 ( .A0(n35598), .A1(n31425), .B0(n16649), .C0(n31424), .Y(
        n15696) );
  INVXL U34540 ( .A(conv_3[6]), .Y(n31429) );
  NAND2XL U34541 ( .A(conv_3[6]), .B(n31427), .Y(n31426) );
  OAI211XL U34542 ( .A0(conv_3[6]), .A1(n31427), .B0(n33157), .C0(n31426), .Y(
        n31428) );
  OAI211XL U34543 ( .A0(n34383), .A1(n31429), .B0(n33468), .C0(n31428), .Y(
        n15742) );
  NAND2XL U34544 ( .A(conv_3[70]), .B(n31433), .Y(n31432) );
  OAI211XL U34545 ( .A0(conv_3[70]), .A1(n31433), .B0(n24499), .C0(n31432), 
        .Y(n31434) );
  OAI211XL U34546 ( .A0(n35598), .A1(n31435), .B0(n33468), .C0(n31434), .Y(
        n15698) );
  NOR2X1 U34547 ( .A(n31437), .B(n31436), .Y(n33797) );
  AOI21XL U34548 ( .A0(n33797), .A1(conv_3[130]), .B0(n35622), .Y(n33709) );
  NOR2X1 U34549 ( .A(n31438), .B(n34783), .Y(n33795) );
  NOR2X1 U34550 ( .A(conv_3[130]), .B(n33795), .Y(n33796) );
  NOR2X1 U34551 ( .A(n33796), .B(n34783), .Y(n33710) );
  NAND2XL U34552 ( .A(conv_3[131]), .B(n31440), .Y(n31439) );
  OAI211XL U34553 ( .A0(conv_3[131]), .A1(n31440), .B0(n16656), .C0(n31439), 
        .Y(n31441) );
  OAI211XL U34554 ( .A0(n35626), .A1(n31442), .B0(n33468), .C0(n31441), .Y(
        n15657) );
  NAND2XL U34555 ( .A(conv_3[305]), .B(n31446), .Y(n31445) );
  OAI211XL U34556 ( .A0(conv_3[305]), .A1(n31446), .B0(n16657), .C0(n31445), 
        .Y(n31447) );
  OAI211XL U34557 ( .A0(n35736), .A1(n31448), .B0(n16649), .C0(n31447), .Y(
        n15543) );
  INVXL U34558 ( .A(conv_3[352]), .Y(n31468) );
  NAND2XL U34559 ( .A(conv_3[351]), .B(n31449), .Y(n31467) );
  AOI21XL U34560 ( .A0(n32130), .A1(n31467), .B0(n31466), .Y(n31452) );
  NAND2XL U34561 ( .A(conv_3[352]), .B(n31452), .Y(n31451) );
  OAI211XL U34562 ( .A0(conv_3[352]), .A1(n31452), .B0(n16656), .C0(n31451), 
        .Y(n31453) );
  OAI211XL U34563 ( .A0(n34746), .A1(n31468), .B0(n16649), .C0(n31453), .Y(
        n15511) );
  AOI21XL U34564 ( .A0(n31455), .A1(n34164), .B0(n31454), .Y(n31457) );
  NAND2XL U34565 ( .A(conv_3[380]), .B(n31457), .Y(n31456) );
  OAI211XL U34566 ( .A0(conv_3[380]), .A1(n31457), .B0(n33788), .C0(n31456), 
        .Y(n31458) );
  OAI211XL U34567 ( .A0(n34168), .A1(n31459), .B0(n16649), .C0(n31458), .Y(
        n15493) );
  AOI21XL U34568 ( .A0(conv_3[384]), .A1(n31502), .B0(n34164), .Y(n31460) );
  AOI21XL U34569 ( .A0(n34164), .A1(n31461), .B0(n31460), .Y(n31463) );
  NAND2XL U34570 ( .A(conv_3[385]), .B(n31463), .Y(n31462) );
  OAI211XL U34571 ( .A0(conv_3[385]), .A1(n31463), .B0(n30090), .C0(n31462), 
        .Y(n31464) );
  OAI211XL U34572 ( .A0(n34168), .A1(n31465), .B0(n33468), .C0(n31464), .Y(
        n15488) );
  NAND2XL U34573 ( .A(conv_3[353]), .B(n33751), .Y(n31486) );
  AOI21XL U34574 ( .A0(conv_3[355]), .A1(n33474), .B0(n33752), .Y(n32129) );
  NAND2XL U34575 ( .A(conv_3[356]), .B(n31470), .Y(n31469) );
  OAI211XL U34576 ( .A0(conv_3[356]), .A1(n31470), .B0(n33712), .C0(n31469), 
        .Y(n31471) );
  OAI211XL U34577 ( .A0(n34746), .A1(n31472), .B0(n33468), .C0(n31471), .Y(
        n15507) );
  OAI21XL U34578 ( .A0(n35599), .A1(n31474), .B0(n31473), .Y(n31476) );
  NAND2XL U34579 ( .A(n31478), .B(n31476), .Y(n31475) );
  OAI211XL U34580 ( .A0(n31478), .A1(n31476), .B0(n33778), .C0(n31475), .Y(
        n31477) );
  OAI211XL U34581 ( .A0(n35598), .A1(n31478), .B0(n16649), .C0(n31477), .Y(
        n15699) );
  NAND2XL U34582 ( .A(conv_3[350]), .B(n31482), .Y(n31481) );
  OAI211XL U34583 ( .A0(conv_3[350]), .A1(n31482), .B0(n33822), .C0(n31481), 
        .Y(n31483) );
  OAI211XL U34584 ( .A0(n34746), .A1(n31484), .B0(n33468), .C0(n31483), .Y(
        n15513) );
  AOI21XL U34585 ( .A0(n32130), .A1(n31486), .B0(n31485), .Y(n31488) );
  NAND2XL U34586 ( .A(conv_3[354]), .B(n31488), .Y(n31487) );
  OAI211XL U34587 ( .A0(conv_3[354]), .A1(n31488), .B0(n32656), .C0(n31487), 
        .Y(n31489) );
  OAI211XL U34588 ( .A0(n34746), .A1(n31490), .B0(n16649), .C0(n31489), .Y(
        n15509) );
  OAI32XL U34589 ( .A0(n32163), .A1(n35600), .A2(conv_3[67]), .B0(n35599), 
        .B1(n31491), .Y(n31493) );
  NAND2XL U34590 ( .A(conv_3[68]), .B(n31493), .Y(n31492) );
  OAI211XL U34591 ( .A0(conv_3[68]), .A1(n31493), .B0(n33157), .C0(n31492), 
        .Y(n31494) );
  OAI211XL U34592 ( .A0(n35598), .A1(n31495), .B0(n33468), .C0(n31494), .Y(
        n15700) );
  INVXL U34593 ( .A(conv_3[309]), .Y(n32540) );
  OAI31XL U34594 ( .A0(conv_3[307]), .A1(conv_3[308]), .A2(n35733), .B0(n35732), .Y(n32535) );
  AOI21XL U34595 ( .A0(conv_3[308]), .A1(n31496), .B0(n35732), .Y(n32536) );
  AOI21XL U34596 ( .A0(n33111), .A1(n35732), .B0(n31497), .Y(n31499) );
  NAND2XL U34597 ( .A(conv_3[312]), .B(n31499), .Y(n31498) );
  OAI211XL U34598 ( .A0(conv_3[312]), .A1(n31499), .B0(n16656), .C0(n31498), 
        .Y(n31500) );
  OAI211XL U34599 ( .A0(n35736), .A1(n33110), .B0(n16649), .C0(n31500), .Y(
        n15536) );
  OAI21XL U34600 ( .A0(n34164), .A1(n31502), .B0(n31501), .Y(n31504) );
  NAND2XL U34601 ( .A(n31506), .B(n31504), .Y(n31503) );
  OAI211XL U34602 ( .A0(n31506), .A1(n31504), .B0(n34028), .C0(n31503), .Y(
        n31505) );
  OAI211XL U34603 ( .A0(n34168), .A1(n31506), .B0(n33468), .C0(n31505), .Y(
        n15489) );
  AOI21XL U34604 ( .A0(n31517), .A1(n31508), .B0(n31507), .Y(n31510) );
  NAND2XL U34605 ( .A(conv_3[456]), .B(n31510), .Y(n31509) );
  OAI211XL U34606 ( .A0(conv_3[456]), .A1(n31510), .B0(n33788), .C0(n31509), 
        .Y(n31511) );
  OAI211XL U34607 ( .A0(n35805), .A1(n31512), .B0(n16649), .C0(n31511), .Y(
        n15442) );
  OAI2BB1XL U34608 ( .A0N(conv_3[460]), .A1N(n31513), .B0(n31517), .Y(n31524)
         );
  AOI32XL U34609 ( .A0(conv_3[461]), .A1(n31517), .A2(n31524), .B0(n33780), 
        .B1(n31519), .Y(n31515) );
  NAND2XL U34610 ( .A(n31518), .B(n31515), .Y(n31514) );
  OAI211XL U34611 ( .A0(n31518), .A1(n31515), .B0(n33822), .C0(n31514), .Y(
        n31516) );
  OAI211XL U34612 ( .A0(n35805), .A1(n31518), .B0(n16649), .C0(n31516), .Y(
        n15436) );
  NAND4XL U34613 ( .A(conv_3[461]), .B(conv_3[462]), .C(n31517), .D(n31524), 
        .Y(n32243) );
  NAND3XL U34614 ( .A(n31519), .B(n33780), .C(n31518), .Y(n32242) );
  NAND2XL U34615 ( .A(n32243), .B(n32242), .Y(n31521) );
  NAND2XL U34616 ( .A(conv_3[463]), .B(n31521), .Y(n31520) );
  OAI211XL U34617 ( .A0(conv_3[463]), .A1(n31521), .B0(n24499), .C0(n31520), 
        .Y(n31522) );
  OAI211XL U34618 ( .A0(n35805), .A1(n32241), .B0(n16649), .C0(n31522), .Y(
        n15435) );
  NAND2XL U34619 ( .A(conv_3[461]), .B(n31526), .Y(n31525) );
  OAI211XL U34620 ( .A0(conv_3[461]), .A1(n31526), .B0(n16657), .C0(n31525), 
        .Y(n31527) );
  OAI211XL U34621 ( .A0(n35805), .A1(n31528), .B0(n16649), .C0(n31527), .Y(
        n15437) );
  NAND2XL U34622 ( .A(conv_3[218]), .B(n32059), .Y(n31537) );
  AOI2BB1XL U34623 ( .A0N(n35660), .A1N(n31542), .B0(n31543), .Y(n31533) );
  NAND2XL U34624 ( .A(conv_3[220]), .B(n31533), .Y(n31532) );
  OAI211XL U34625 ( .A0(conv_3[220]), .A1(n31533), .B0(n33912), .C0(n31532), 
        .Y(n31534) );
  OAI211XL U34626 ( .A0(n35665), .A1(n31535), .B0(n33468), .C0(n31534), .Y(
        n15598) );
  AOI21XL U34627 ( .A0(n34649), .A1(n31537), .B0(n31536), .Y(n31539) );
  NAND2XL U34628 ( .A(conv_3[219]), .B(n31539), .Y(n31538) );
  OAI211XL U34629 ( .A0(conv_3[219]), .A1(n31539), .B0(n33912), .C0(n31538), 
        .Y(n31540) );
  OAI211XL U34630 ( .A0(n35665), .A1(n31541), .B0(n33468), .C0(n31540), .Y(
        n15599) );
  OAI2BB1XL U34631 ( .A0N(conv_3[220]), .A1N(n31542), .B0(n34649), .Y(n35667)
         );
  NAND4XL U34632 ( .A(conv_3[221]), .B(conv_3[222]), .C(n34649), .D(n35667), 
        .Y(n32138) );
  OAI21XL U34633 ( .A0(conv_3[220]), .A1(n31543), .B0(n35660), .Y(n35666) );
  NAND3XL U34634 ( .A(n35668), .B(n35660), .C(n34653), .Y(n32137) );
  NAND2XL U34635 ( .A(n32138), .B(n32137), .Y(n31545) );
  NAND2XL U34636 ( .A(conv_3[223]), .B(n31545), .Y(n31544) );
  OAI211XL U34637 ( .A0(conv_3[223]), .A1(n31545), .B0(n33912), .C0(n31544), 
        .Y(n31546) );
  OAI211XL U34638 ( .A0(n35665), .A1(n32136), .B0(n33468), .C0(n31546), .Y(
        n15595) );
  INVXL U34639 ( .A(conv_3[491]), .Y(n31554) );
  OAI21XL U34640 ( .A0(conv_3[490]), .A1(n35829), .B0(n35831), .Y(n31553) );
  OAI2BB1XL U34641 ( .A0N(conv_3[490]), .A1N(n35830), .B0(n35823), .Y(n32227)
         );
  NAND2XL U34642 ( .A(n31553), .B(n32227), .Y(n31551) );
  NAND2XL U34643 ( .A(n31554), .B(n31551), .Y(n31550) );
  OAI211XL U34644 ( .A0(n31554), .A1(n31551), .B0(n32181), .C0(n31550), .Y(
        n31552) );
  OAI211XL U34645 ( .A0(n35826), .A1(n31554), .B0(n16649), .C0(n31552), .Y(
        n15417) );
  INVXL U34646 ( .A(conv_3[492]), .Y(n32229) );
  NAND2XL U34647 ( .A(n31554), .B(n31553), .Y(n31555) );
  NAND2XL U34648 ( .A(n35831), .B(n31555), .Y(n32228) );
  AOI32XL U34649 ( .A0(conv_3[491]), .A1(n32228), .A2(n32227), .B0(n35831), 
        .B1(n32228), .Y(n31557) );
  NAND2XL U34650 ( .A(n32229), .B(n31557), .Y(n31556) );
  OAI211XL U34651 ( .A0(n32229), .A1(n31557), .B0(n16656), .C0(n31556), .Y(
        n31558) );
  OAI211XL U34652 ( .A0(n35826), .A1(n32229), .B0(n16649), .C0(n31558), .Y(
        n15416) );
  AOI2BB1XL U34653 ( .A0N(n35639), .A1N(n31567), .B0(n31568), .Y(n31564) );
  NAND2XL U34654 ( .A(conv_3[171]), .B(n31564), .Y(n31563) );
  OAI211XL U34655 ( .A0(conv_3[171]), .A1(n31564), .B0(n30090), .C0(n31563), 
        .Y(n31565) );
  OAI211XL U34656 ( .A0(n35630), .A1(n31566), .B0(n33468), .C0(n31565), .Y(
        n15632) );
  INVXL U34657 ( .A(conv_3[176]), .Y(n31572) );
  OAI2BB1XL U34658 ( .A0N(n31567), .A1N(conv_3[171]), .B0(n32221), .Y(n35631)
         );
  OAI21XL U34659 ( .A0(conv_3[171]), .A1(n31568), .B0(n35639), .Y(n35629) );
  NOR2BX1 U34660 ( .AN(n35629), .B(conv_3[172]), .Y(n35632) );
  AOI31XL U34661 ( .A0(conv_3[175]), .A1(conv_3[174]), .A2(n31573), .B0(n35639), .Y(n31578) );
  NAND2XL U34662 ( .A(conv_3[176]), .B(n31570), .Y(n31569) );
  OAI211XL U34663 ( .A0(conv_3[176]), .A1(n31570), .B0(n33982), .C0(n31569), 
        .Y(n31571) );
  OAI211XL U34664 ( .A0(n35630), .A1(n31572), .B0(n33468), .C0(n31571), .Y(
        n15627) );
  INVXL U34665 ( .A(conv_3[174]), .Y(n35635) );
  AOI21XL U34666 ( .A0(n31573), .A1(n35639), .B0(n35636), .Y(n31575) );
  NAND2XL U34667 ( .A(conv_3[174]), .B(n31575), .Y(n31574) );
  OAI211XL U34668 ( .A0(conv_3[174]), .A1(n31575), .B0(n34028), .C0(n31574), 
        .Y(n31576) );
  OAI211XL U34669 ( .A0(n35630), .A1(n35635), .B0(n33468), .C0(n31576), .Y(
        n15629) );
  AOI2BB1XL U34670 ( .A0N(n35639), .A1N(n32220), .B0(n32222), .Y(n31581) );
  NAND2XL U34671 ( .A(conv_3[177]), .B(n31581), .Y(n31580) );
  OAI211XL U34672 ( .A0(conv_3[177]), .A1(n31581), .B0(n33788), .C0(n31580), 
        .Y(n31582) );
  OAI211XL U34673 ( .A0(n35630), .A1(n31583), .B0(n33468), .C0(n31582), .Y(
        n15626) );
  NAND2XL U34674 ( .A(conv_3[170]), .B(n31587), .Y(n31586) );
  OAI211XL U34675 ( .A0(conv_3[170]), .A1(n31587), .B0(n34028), .C0(n31586), 
        .Y(n31588) );
  OAI211XL U34676 ( .A0(n35630), .A1(n31589), .B0(n33468), .C0(n31588), .Y(
        n15633) );
  OAI21XL U34677 ( .A0(n31597), .A1(conv_3[187]), .B0(n32649), .Y(n31590) );
  OAI21XL U34678 ( .A0(n32649), .A1(n31591), .B0(n31590), .Y(n31593) );
  NAND2XL U34679 ( .A(n31595), .B(n31593), .Y(n31592) );
  OAI211XL U34680 ( .A0(n31595), .A1(n31593), .B0(n33982), .C0(n31592), .Y(
        n31594) );
  OAI211XL U34681 ( .A0(n34704), .A1(n31595), .B0(n33468), .C0(n31594), .Y(
        n15620) );
  AOI21XL U34682 ( .A0(n31597), .A1(n32649), .B0(n31596), .Y(n31599) );
  NAND2XL U34683 ( .A(conv_3[187]), .B(n31599), .Y(n31598) );
  OAI211XL U34684 ( .A0(conv_3[187]), .A1(n31599), .B0(n34028), .C0(n31598), 
        .Y(n31600) );
  OAI211XL U34685 ( .A0(n34704), .A1(n31601), .B0(n33468), .C0(n31600), .Y(
        n15621) );
  NAND2XL U34686 ( .A(conv_3[191]), .B(n31604), .Y(n31603) );
  OAI211XL U34687 ( .A0(conv_3[191]), .A1(n31604), .B0(n33982), .C0(n31603), 
        .Y(n31605) );
  OAI211XL U34688 ( .A0(n34704), .A1(n31606), .B0(n33468), .C0(n31605), .Y(
        n15617) );
  OAI32XL U34689 ( .A0(n32649), .A1(n31609), .A2(n31608), .B0(n32207), .B1(
        n31607), .Y(n31611) );
  NAND2XL U34690 ( .A(conv_3[190]), .B(n31611), .Y(n31610) );
  OAI211XL U34691 ( .A0(conv_3[190]), .A1(n31611), .B0(n33788), .C0(n31610), 
        .Y(n31612) );
  OAI211XL U34692 ( .A0(n34704), .A1(n31613), .B0(n33468), .C0(n31612), .Y(
        n15618) );
  NAND2XL U34693 ( .A(conv_3[185]), .B(n31617), .Y(n31616) );
  OAI211XL U34694 ( .A0(conv_3[185]), .A1(n31617), .B0(n33982), .C0(n31616), 
        .Y(n31618) );
  OAI211XL U34695 ( .A0(n34704), .A1(n31619), .B0(n33468), .C0(n31618), .Y(
        n15623) );
  INVXL U34696 ( .A(conv_3[193]), .Y(n32205) );
  NAND2XL U34697 ( .A(n32208), .B(n32207), .Y(n32206) );
  OAI21XL U34698 ( .A0(n32208), .A1(n32207), .B0(n32206), .Y(n31623) );
  NAND2XL U34699 ( .A(conv_3[193]), .B(n31623), .Y(n31622) );
  OAI211XL U34700 ( .A0(conv_3[193]), .A1(n31623), .B0(n32181), .C0(n31622), 
        .Y(n31624) );
  OAI211XL U34701 ( .A0(n34704), .A1(n32205), .B0(n33468), .C0(n31624), .Y(
        n15615) );
  INVXL U34702 ( .A(conv_3[367]), .Y(n31659) );
  NAND2XL U34703 ( .A(conv_3[366]), .B(n31661), .Y(n31655) );
  NAND2XL U34704 ( .A(conv_3[368]), .B(n31649), .Y(n35760) );
  OAI2BB1XL U34705 ( .A0N(conv_3[370]), .A1N(n33832), .B0(n35761), .Y(n31642)
         );
  AOI32XL U34706 ( .A0(conv_3[371]), .A1(n35761), .A2(n31642), .B0(n33833), 
        .B1(n31644), .Y(n31629) );
  NAND2XL U34707 ( .A(n31643), .B(n31629), .Y(n31628) );
  OAI211XL U34708 ( .A0(n31643), .A1(n31629), .B0(n30090), .C0(n31628), .Y(
        n31630) );
  OAI211XL U34709 ( .A0(n35764), .A1(n31643), .B0(n33468), .C0(n31630), .Y(
        n15496) );
  NAND2XL U34710 ( .A(conv_3[371]), .B(n31633), .Y(n31632) );
  OAI211XL U34711 ( .A0(conv_3[371]), .A1(n31633), .B0(n33778), .C0(n31632), 
        .Y(n31634) );
  OAI211XL U34712 ( .A0(n35764), .A1(n31635), .B0(n16649), .C0(n31634), .Y(
        n15497) );
  NAND2XL U34713 ( .A(conv_3[365]), .B(n31639), .Y(n31638) );
  OAI211XL U34714 ( .A0(conv_3[365]), .A1(n31639), .B0(n16657), .C0(n31638), 
        .Y(n31640) );
  OAI211XL U34715 ( .A0(n35764), .A1(n31641), .B0(n33468), .C0(n31640), .Y(
        n15503) );
  NAND4XL U34716 ( .A(conv_3[371]), .B(conv_3[372]), .C(n35761), .D(n31642), 
        .Y(n32123) );
  NAND3XL U34717 ( .A(n31644), .B(n33833), .C(n31643), .Y(n32122) );
  NAND2XL U34718 ( .A(n32123), .B(n32122), .Y(n31646) );
  NAND2XL U34719 ( .A(conv_3[373]), .B(n31646), .Y(n31645) );
  OAI211XL U34720 ( .A0(conv_3[373]), .A1(n31646), .B0(n33982), .C0(n31645), 
        .Y(n31647) );
  OAI211XL U34721 ( .A0(n35764), .A1(n32121), .B0(n16649), .C0(n31647), .Y(
        n15495) );
  INVXL U34722 ( .A(conv_3[368]), .Y(n31653) );
  AOI2BB1XL U34723 ( .A0N(n33833), .A1N(n31649), .B0(n31648), .Y(n31651) );
  NAND2XL U34724 ( .A(conv_3[368]), .B(n31651), .Y(n31650) );
  OAI211XL U34725 ( .A0(conv_3[368]), .A1(n31651), .B0(n33157), .C0(n31650), 
        .Y(n31652) );
  OAI211XL U34726 ( .A0(n35764), .A1(n31653), .B0(n16649), .C0(n31652), .Y(
        n15500) );
  AOI21XL U34727 ( .A0(n35761), .A1(n31655), .B0(n31654), .Y(n31657) );
  NAND2XL U34728 ( .A(conv_3[367]), .B(n31657), .Y(n31656) );
  OAI211XL U34729 ( .A0(conv_3[367]), .A1(n31657), .B0(n33788), .C0(n31656), 
        .Y(n31658) );
  OAI211XL U34730 ( .A0(n35764), .A1(n31659), .B0(n33468), .C0(n31658), .Y(
        n15501) );
  INVXL U34731 ( .A(conv_3[366]), .Y(n31665) );
  AOI2BB1XL U34732 ( .A0N(n33833), .A1N(n31661), .B0(n31660), .Y(n31663) );
  NAND2XL U34733 ( .A(conv_3[366]), .B(n31663), .Y(n31662) );
  OAI211XL U34734 ( .A0(conv_3[366]), .A1(n31663), .B0(n32611), .C0(n31662), 
        .Y(n31664) );
  OAI211XL U34735 ( .A0(n35764), .A1(n31665), .B0(n33468), .C0(n31664), .Y(
        n15502) );
  INVXL U34736 ( .A(conv_3[99]), .Y(n35617) );
  NAND2XL U34737 ( .A(conv_3[96]), .B(n33743), .Y(n31674) );
  NAND2XL U34738 ( .A(conv_3[98]), .B(n31686), .Y(n35614) );
  NAND2XL U34739 ( .A(conv_3[100]), .B(n31670), .Y(n31669) );
  OAI211XL U34740 ( .A0(conv_3[100]), .A1(n31670), .B0(n16656), .C0(n31669), 
        .Y(n31671) );
  OAI211XL U34741 ( .A0(n35618), .A1(n31672), .B0(n16649), .C0(n31671), .Y(
        n15678) );
  AOI21XL U34742 ( .A0(n35615), .A1(n31674), .B0(n31673), .Y(n31676) );
  NAND2XL U34743 ( .A(conv_3[97]), .B(n31676), .Y(n31675) );
  OAI211XL U34744 ( .A0(conv_3[97]), .A1(n31676), .B0(n33912), .C0(n31675), 
        .Y(n31677) );
  OAI211XL U34745 ( .A0(n35618), .A1(n31678), .B0(n33468), .C0(n31677), .Y(
        n15681) );
  NAND2XL U34746 ( .A(conv_3[95]), .B(n31682), .Y(n31681) );
  OAI211XL U34747 ( .A0(conv_3[95]), .A1(n31682), .B0(n33778), .C0(n31681), 
        .Y(n31683) );
  OAI211XL U34748 ( .A0(n35618), .A1(n31684), .B0(n33468), .C0(n31683), .Y(
        n15683) );
  INVXL U34749 ( .A(conv_3[98]), .Y(n31690) );
  AOI2BB1XL U34750 ( .A0N(n34186), .A1N(n31686), .B0(n31685), .Y(n31688) );
  NAND2XL U34751 ( .A(conv_3[98]), .B(n31688), .Y(n31687) );
  OAI211XL U34752 ( .A0(conv_3[98]), .A1(n31688), .B0(n16657), .C0(n31687), 
        .Y(n31689) );
  OAI211XL U34753 ( .A0(n35618), .A1(n31690), .B0(n16649), .C0(n31689), .Y(
        n15680) );
  INVXL U34754 ( .A(conv_3[430]), .Y(n31700) );
  INVXL U34755 ( .A(conv_3[427]), .Y(n35770) );
  NAND2XL U34756 ( .A(conv_3[426]), .B(n33789), .Y(n35768) );
  NAND2XL U34757 ( .A(conv_3[428]), .B(n31702), .Y(n35774) );
  AOI2BB1XL U34758 ( .A0N(n33790), .A1N(n31725), .B0(n31726), .Y(n31698) );
  NAND2XL U34759 ( .A(conv_3[430]), .B(n31698), .Y(n31697) );
  OAI211XL U34760 ( .A0(conv_3[430]), .A1(n31698), .B0(n33788), .C0(n31697), 
        .Y(n31699) );
  OAI211XL U34761 ( .A0(n35778), .A1(n31700), .B0(n16649), .C0(n31699), .Y(
        n15458) );
  AOI2BB1XL U34762 ( .A0N(n33790), .A1N(n31702), .B0(n31701), .Y(n31704) );
  NAND2XL U34763 ( .A(conv_3[428]), .B(n31704), .Y(n31703) );
  OAI211XL U34764 ( .A0(conv_3[428]), .A1(n31704), .B0(n34666), .C0(n31703), 
        .Y(n31705) );
  OAI211XL U34765 ( .A0(n35778), .A1(n31706), .B0(n16649), .C0(n31705), .Y(
        n15460) );
  AOI21XL U34766 ( .A0(n32789), .A1(n31708), .B0(n31707), .Y(n31710) );
  NAND2XL U34767 ( .A(conv_3[144]), .B(n31710), .Y(n31709) );
  OAI211XL U34768 ( .A0(conv_3[144]), .A1(n31710), .B0(n34028), .C0(n31709), 
        .Y(n31711) );
  OAI211XL U34769 ( .A0(n34737), .A1(n31712), .B0(n33468), .C0(n31711), .Y(
        n15649) );
  NAND2XL U34770 ( .A(conv_3[141]), .B(n31716), .Y(n31715) );
  OAI211XL U34771 ( .A0(conv_3[141]), .A1(n31716), .B0(n32181), .C0(n31715), 
        .Y(n31717) );
  OAI211XL U34772 ( .A0(n34737), .A1(n31718), .B0(n16649), .C0(n31717), .Y(
        n15652) );
  INVXL U34773 ( .A(conv_3[143]), .Y(n31724) );
  AOI21XL U34774 ( .A0(n31720), .A1(n33466), .B0(n31719), .Y(n31722) );
  NAND2XL U34775 ( .A(conv_3[143]), .B(n31722), .Y(n31721) );
  OAI211XL U34776 ( .A0(conv_3[143]), .A1(n31722), .B0(n34028), .C0(n31721), 
        .Y(n31723) );
  OAI211XL U34777 ( .A0(n34737), .A1(n31724), .B0(n33468), .C0(n31723), .Y(
        n15650) );
  OAI2BB1XL U34778 ( .A0N(conv_3[430]), .A1N(n31725), .B0(n35775), .Y(n32582)
         );
  NAND2XL U34779 ( .A(conv_3[431]), .B(n31728), .Y(n31727) );
  OAI211XL U34780 ( .A0(conv_3[431]), .A1(n31728), .B0(n33788), .C0(n31727), 
        .Y(n31729) );
  OAI211XL U34781 ( .A0(n35778), .A1(n31730), .B0(n16649), .C0(n31729), .Y(
        n15457) );
  INVXL U34782 ( .A(conv_3[283]), .Y(n32257) );
  AOI21XL U34783 ( .A0(n31732), .A1(n31731), .B0(n32599), .Y(n31744) );
  NAND2XL U34784 ( .A(conv_3[275]), .B(n31733), .Y(n31745) );
  INVXL U34785 ( .A(conv_3[276]), .Y(n31749) );
  AOI21XL U34786 ( .A0(n31751), .A1(conv_3[277]), .B0(n32618), .Y(n31739) );
  OAI2BB1XL U34787 ( .A0N(conv_3[280]), .A1N(n31757), .B0(n32599), .Y(n32598)
         );
  NAND4XL U34788 ( .A(conv_3[281]), .B(conv_3[282]), .C(n32599), .D(n32598), 
        .Y(n32259) );
  NAND3XL U34789 ( .A(n32597), .B(n32618), .C(n32603), .Y(n32258) );
  NAND2XL U34790 ( .A(n32259), .B(n32258), .Y(n31736) );
  NAND2XL U34791 ( .A(conv_3[283]), .B(n31736), .Y(n31734) );
  OAI211XL U34792 ( .A0(conv_3[283]), .A1(n31736), .B0(n31735), .C0(n31734), 
        .Y(n31737) );
  OAI211XL U34793 ( .A0(n34709), .A1(n32257), .B0(n33468), .C0(n31737), .Y(
        n15555) );
  NAND2XL U34794 ( .A(conv_3[278]), .B(n31741), .Y(n31740) );
  OAI211XL U34795 ( .A0(conv_3[278]), .A1(n31741), .B0(n32611), .C0(n31740), 
        .Y(n31742) );
  OAI211XL U34796 ( .A0(n34709), .A1(n31743), .B0(n33468), .C0(n31742), .Y(
        n15560) );
  AOI21XL U34797 ( .A0(n32599), .A1(n31745), .B0(n31744), .Y(n31747) );
  NAND2XL U34798 ( .A(conv_3[276]), .B(n31747), .Y(n31746) );
  OAI211XL U34799 ( .A0(conv_3[276]), .A1(n31747), .B0(n33982), .C0(n31746), 
        .Y(n31748) );
  OAI211XL U34800 ( .A0(n34709), .A1(n31749), .B0(n16649), .C0(n31748), .Y(
        n15562) );
  INVXL U34801 ( .A(conv_3[277]), .Y(n31755) );
  AOI2BB1XL U34802 ( .A0N(n32618), .A1N(n31751), .B0(n31750), .Y(n31753) );
  NAND2XL U34803 ( .A(conv_3[277]), .B(n31753), .Y(n31752) );
  OAI211XL U34804 ( .A0(conv_3[277]), .A1(n31753), .B0(n33982), .C0(n31752), 
        .Y(n31754) );
  OAI211XL U34805 ( .A0(n34709), .A1(n31755), .B0(n33468), .C0(n31754), .Y(
        n15561) );
  INVXL U34806 ( .A(conv_3[280]), .Y(n31761) );
  AOI21XL U34807 ( .A0(n31757), .A1(n32618), .B0(n31756), .Y(n31759) );
  NAND2XL U34808 ( .A(conv_3[280]), .B(n31759), .Y(n31758) );
  OAI211XL U34809 ( .A0(conv_3[280]), .A1(n31759), .B0(n16657), .C0(n31758), 
        .Y(n31760) );
  OAI211XL U34810 ( .A0(n34709), .A1(n31761), .B0(n16649), .C0(n31760), .Y(
        n15558) );
  INVXL U34811 ( .A(conv_3[281]), .Y(n31766) );
  NOR2BXL U34812 ( .AN(n32598), .B(n31762), .Y(n31764) );
  NAND2XL U34813 ( .A(conv_3[281]), .B(n31764), .Y(n31763) );
  OAI211XL U34814 ( .A0(conv_3[281]), .A1(n31764), .B0(n32181), .C0(n31763), 
        .Y(n31765) );
  OAI211XL U34815 ( .A0(n34709), .A1(n31766), .B0(n16649), .C0(n31765), .Y(
        n15557) );
  NAND2XL U34816 ( .A(n31786), .B(n31769), .Y(n31775) );
  NOR2BXL U34817 ( .AN(n31775), .B(n31774), .Y(n31771) );
  NAND2XL U34818 ( .A(conv_3[110]), .B(n31771), .Y(n31770) );
  OAI211XL U34819 ( .A0(conv_3[110]), .A1(n31771), .B0(n32611), .C0(n31770), 
        .Y(n31772) );
  OAI211XL U34820 ( .A0(n34200), .A1(n31773), .B0(n16649), .C0(n31772), .Y(
        n15673) );
  INVXL U34821 ( .A(conv_3[116]), .Y(n31779) );
  NAND2XL U34822 ( .A(conv_3[110]), .B(n31775), .Y(n31785) );
  INVXL U34823 ( .A(conv_3[111]), .Y(n31790) );
  AOI21XL U34824 ( .A0(conv_3[115]), .A1(n32636), .B0(n34196), .Y(n31780) );
  AOI221XL U34825 ( .A0(conv_3[115]), .A1(n34196), .B0(n32636), .B1(n34196), 
        .C0(n31780), .Y(n31777) );
  NAND2XL U34826 ( .A(conv_3[116]), .B(n31777), .Y(n31776) );
  OAI211XL U34827 ( .A0(conv_3[116]), .A1(n31777), .B0(n33157), .C0(n31776), 
        .Y(n31778) );
  OAI211XL U34828 ( .A0(n34200), .A1(n31779), .B0(n16649), .C0(n31778), .Y(
        n15667) );
  INVXL U34829 ( .A(conv_3[118]), .Y(n32264) );
  NAND3XL U34830 ( .A(conv_3[117]), .B(n34195), .C(n31786), .Y(n32266) );
  OAI31XL U34831 ( .A0(conv_3[116]), .A1(conv_3[115]), .A2(n32636), .B0(n34196), .Y(n34194) );
  NAND3XL U34832 ( .A(n34196), .B(n34201), .C(n34194), .Y(n32265) );
  NAND2XL U34833 ( .A(n32266), .B(n32265), .Y(n31782) );
  NAND2XL U34834 ( .A(conv_3[118]), .B(n31782), .Y(n31781) );
  OAI211XL U34835 ( .A0(conv_3[118]), .A1(n31782), .B0(n30090), .C0(n31781), 
        .Y(n31783) );
  OAI211XL U34836 ( .A0(n34200), .A1(n32264), .B0(n33468), .C0(n31783), .Y(
        n15665) );
  AOI21XL U34837 ( .A0(n31786), .A1(n31785), .B0(n31784), .Y(n31788) );
  NAND2XL U34838 ( .A(conv_3[111]), .B(n31788), .Y(n31787) );
  OAI211XL U34839 ( .A0(conv_3[111]), .A1(n31788), .B0(n33778), .C0(n31787), 
        .Y(n31789) );
  OAI211XL U34840 ( .A0(n34200), .A1(n31790), .B0(n16649), .C0(n31789), .Y(
        n15672) );
  INVXL U34841 ( .A(conv_3[113]), .Y(n31796) );
  NAND2XL U34842 ( .A(conv_3[113]), .B(n31794), .Y(n31793) );
  OAI211XL U34843 ( .A0(conv_3[113]), .A1(n31794), .B0(n33788), .C0(n31793), 
        .Y(n31795) );
  OAI211XL U34844 ( .A0(n34200), .A1(n31796), .B0(n33468), .C0(n31795), .Y(
        n15670) );
  AOI2BB1XL U34845 ( .A0N(n34196), .A1N(n31798), .B0(n31797), .Y(n31800) );
  NAND2XL U34846 ( .A(conv_3[112]), .B(n31800), .Y(n31799) );
  OAI211XL U34847 ( .A0(conv_3[112]), .A1(n31800), .B0(n33982), .C0(n31799), 
        .Y(n31801) );
  OAI211XL U34848 ( .A0(n34200), .A1(n31802), .B0(n33468), .C0(n31801), .Y(
        n15671) );
  INVXL U34849 ( .A(conv_3[80]), .Y(n34154) );
  NAND2XL U34850 ( .A(conv_3[81]), .B(n31822), .Y(n31834) );
  NAND2XL U34851 ( .A(conv_3[83]), .B(n31811), .Y(n35606) );
  AOI2BB1XL U34852 ( .A0N(n31842), .A1N(n31817), .B0(n31816), .Y(n31807) );
  NAND2XL U34853 ( .A(conv_3[85]), .B(n31807), .Y(n31806) );
  OAI211XL U34854 ( .A0(conv_3[85]), .A1(n31807), .B0(n32660), .C0(n31806), 
        .Y(n31808) );
  OAI211XL U34855 ( .A0(n35610), .A1(n31809), .B0(n16649), .C0(n31808), .Y(
        n15688) );
  INVXL U34856 ( .A(conv_3[83]), .Y(n31815) );
  AOI2BB1XL U34857 ( .A0N(n31842), .A1N(n31811), .B0(n31810), .Y(n31813) );
  NAND2XL U34858 ( .A(conv_3[83]), .B(n31813), .Y(n31812) );
  OAI211XL U34859 ( .A0(conv_3[83]), .A1(n31813), .B0(n30090), .C0(n31812), 
        .Y(n31814) );
  OAI211XL U34860 ( .A0(n35610), .A1(n31815), .B0(n16649), .C0(n31814), .Y(
        n15690) );
  INVXL U34861 ( .A(conv_3[86]), .Y(n31828) );
  OAI21XL U34862 ( .A0(conv_3[85]), .A1(n31816), .B0(n31842), .Y(n31827) );
  OAI2BB1XL U34863 ( .A0N(conv_3[85]), .A1N(n31817), .B0(n35607), .Y(n31839)
         );
  NAND2XL U34864 ( .A(n31827), .B(n31839), .Y(n31819) );
  NAND2XL U34865 ( .A(n31828), .B(n31819), .Y(n31818) );
  OAI211XL U34866 ( .A0(n31828), .A1(n31819), .B0(n32181), .C0(n31818), .Y(
        n31820) );
  OAI211XL U34867 ( .A0(n35610), .A1(n31828), .B0(n33468), .C0(n31820), .Y(
        n15687) );
  INVXL U34868 ( .A(conv_3[81]), .Y(n31826) );
  AOI2BB1XL U34869 ( .A0N(n31842), .A1N(n31822), .B0(n31821), .Y(n31824) );
  NAND2XL U34870 ( .A(conv_3[81]), .B(n31824), .Y(n31823) );
  OAI211XL U34871 ( .A0(conv_3[81]), .A1(n31824), .B0(n16657), .C0(n31823), 
        .Y(n31825) );
  OAI211XL U34872 ( .A0(n35610), .A1(n31826), .B0(n16649), .C0(n31825), .Y(
        n15692) );
  INVXL U34873 ( .A(conv_3[87]), .Y(n31841) );
  NAND2XL U34874 ( .A(n31828), .B(n31827), .Y(n31829) );
  AOI32XL U34875 ( .A0(conv_3[86]), .A1(n31840), .A2(n31839), .B0(n31842), 
        .B1(n31840), .Y(n31831) );
  NAND2XL U34876 ( .A(n31841), .B(n31831), .Y(n31830) );
  OAI211XL U34877 ( .A0(n31841), .A1(n31831), .B0(n33712), .C0(n31830), .Y(
        n31832) );
  OAI211XL U34878 ( .A0(n35610), .A1(n31841), .B0(n16649), .C0(n31832), .Y(
        n15686) );
  AOI21XL U34879 ( .A0(n35607), .A1(n31834), .B0(n31833), .Y(n31836) );
  NAND2XL U34880 ( .A(conv_3[82]), .B(n31836), .Y(n31835) );
  OAI211XL U34881 ( .A0(conv_3[82]), .A1(n31836), .B0(n32656), .C0(n31835), 
        .Y(n31837) );
  OAI211XL U34882 ( .A0(n35610), .A1(n31838), .B0(n33468), .C0(n31837), .Y(
        n15691) );
  NAND4XL U34883 ( .A(conv_3[86]), .B(conv_3[87]), .C(n35607), .D(n31839), .Y(
        n32152) );
  NAND3XL U34884 ( .A(n31842), .B(n31841), .C(n31840), .Y(n32151) );
  NAND2XL U34885 ( .A(n32152), .B(n32151), .Y(n31844) );
  NAND2XL U34886 ( .A(conv_3[88]), .B(n31844), .Y(n31843) );
  OAI211XL U34887 ( .A0(conv_3[88]), .A1(n31844), .B0(n28751), .C0(n31843), 
        .Y(n31845) );
  OAI211XL U34888 ( .A0(n35610), .A1(n32150), .B0(n33468), .C0(n31845), .Y(
        n15685) );
  INVXL U34889 ( .A(conv_3[208]), .Y(n32271) );
  OAI2BB1XL U34890 ( .A0N(conv_3[205]), .A1N(n35652), .B0(n31848), .Y(n31859)
         );
  NAND4XL U34891 ( .A(conv_3[206]), .B(conv_3[207]), .C(n31848), .D(n31859), 
        .Y(n32273) );
  OAI21XL U34892 ( .A0(conv_3[205]), .A1(n35651), .B0(n35653), .Y(n31854) );
  NAND2XL U34893 ( .A(n31858), .B(n31854), .Y(n31850) );
  NAND3XL U34894 ( .A(n35653), .B(n31864), .C(n31860), .Y(n32272) );
  NAND2XL U34895 ( .A(n32273), .B(n32272), .Y(n31852) );
  NAND2XL U34896 ( .A(conv_3[208]), .B(n31852), .Y(n31851) );
  OAI211XL U34897 ( .A0(conv_3[208]), .A1(n31852), .B0(n33912), .C0(n31851), 
        .Y(n31853) );
  OAI211XL U34898 ( .A0(n35646), .A1(n32271), .B0(n33468), .C0(n31853), .Y(
        n15605) );
  NAND2XL U34899 ( .A(n31854), .B(n31859), .Y(n31856) );
  NAND2XL U34900 ( .A(n31858), .B(n31856), .Y(n31855) );
  OAI211XL U34901 ( .A0(n31858), .A1(n31856), .B0(n31735), .C0(n31855), .Y(
        n31857) );
  OAI211XL U34902 ( .A0(n35646), .A1(n31858), .B0(n33468), .C0(n31857), .Y(
        n15607) );
  AOI32XL U34903 ( .A0(conv_3[206]), .A1(n31860), .A2(n31859), .B0(n35653), 
        .B1(n31860), .Y(n31862) );
  NAND2XL U34904 ( .A(n31864), .B(n31862), .Y(n31861) );
  OAI211XL U34905 ( .A0(n31864), .A1(n31862), .B0(n33912), .C0(n31861), .Y(
        n31863) );
  OAI211XL U34906 ( .A0(n35646), .A1(n31864), .B0(n33468), .C0(n31863), .Y(
        n15606) );
  INVXL U34907 ( .A(conv_3[201]), .Y(n31870) );
  NAND2XL U34908 ( .A(conv_3[201]), .B(n31868), .Y(n31867) );
  OAI211XL U34909 ( .A0(conv_3[201]), .A1(n31868), .B0(n24499), .C0(n31867), 
        .Y(n31869) );
  OAI211XL U34910 ( .A0(n35646), .A1(n31870), .B0(n33468), .C0(n31869), .Y(
        n15612) );
  INVXL U34911 ( .A(conv_3[298]), .Y(n32234) );
  NAND2XL U34912 ( .A(n31890), .B(conv_3[291]), .Y(n31883) );
  INVXL U34913 ( .A(conv_3[292]), .Y(n31887) );
  INVXL U34914 ( .A(n35720), .Y(n31896) );
  OAI31XL U34915 ( .A0(conv_3[290]), .A1(n31888), .A2(conv_3[291]), .B0(n35720), .Y(n31882) );
  AOI21XL U34916 ( .A0(n31887), .A1(n31882), .B0(n31896), .Y(n35718) );
  OAI21XL U34917 ( .A0(conv_3[293]), .A1(n35718), .B0(n35720), .Y(n35725) );
  NAND4XL U34918 ( .A(conv_3[297]), .B(conv_3[296]), .C(n34479), .D(n31896), 
        .Y(n32236) );
  NAND2XL U34919 ( .A(n32236), .B(n32235), .Y(n31875) );
  NAND2XL U34920 ( .A(conv_3[298]), .B(n31875), .Y(n31874) );
  OAI211XL U34921 ( .A0(conv_3[298]), .A1(n31875), .B0(n34666), .C0(n31874), 
        .Y(n31876) );
  OAI211XL U34922 ( .A0(n35726), .A1(n32234), .B0(n16649), .C0(n31876), .Y(
        n15545) );
  AOI21XL U34923 ( .A0(n31888), .A1(n35720), .B0(n31877), .Y(n31879) );
  NAND2XL U34924 ( .A(conv_3[290]), .B(n31879), .Y(n31878) );
  OAI211XL U34925 ( .A0(conv_3[290]), .A1(n31879), .B0(n16656), .C0(n31878), 
        .Y(n31880) );
  OAI211XL U34926 ( .A0(n35726), .A1(n31881), .B0(n33468), .C0(n31880), .Y(
        n15553) );
  OAI2BB1XL U34927 ( .A0N(n31896), .A1N(n31883), .B0(n31882), .Y(n31885) );
  NAND2XL U34928 ( .A(n31887), .B(n31885), .Y(n31884) );
  OAI211XL U34929 ( .A0(n31887), .A1(n31885), .B0(n34666), .C0(n31884), .Y(
        n31886) );
  OAI211XL U34930 ( .A0(n35726), .A1(n31887), .B0(n33468), .C0(n31886), .Y(
        n15551) );
  INVXL U34931 ( .A(conv_3[291]), .Y(n31894) );
  AOI2BB1XL U34932 ( .A0N(n31888), .A1N(conv_3[290]), .B0(n31896), .Y(n31889)
         );
  AOI2BB1XL U34933 ( .A0N(n35720), .A1N(n31890), .B0(n31889), .Y(n31892) );
  NAND2XL U34934 ( .A(conv_3[291]), .B(n31892), .Y(n31891) );
  OAI211XL U34935 ( .A0(conv_3[291]), .A1(n31892), .B0(n34666), .C0(n31891), 
        .Y(n31893) );
  OAI211XL U34936 ( .A0(n35726), .A1(n31894), .B0(n16649), .C0(n31893), .Y(
        n15552) );
  INVXL U34937 ( .A(conv_3[297]), .Y(n31900) );
  NAND2XL U34938 ( .A(n34479), .B(conv_3[296]), .Y(n31895) );
  OAI32XL U34939 ( .A0(n31896), .A1(n34479), .A2(conv_3[296]), .B0(n35720), 
        .B1(n31895), .Y(n31898) );
  NAND2XL U34940 ( .A(conv_3[297]), .B(n31898), .Y(n31897) );
  OAI211XL U34941 ( .A0(conv_3[297]), .A1(n31898), .B0(n34666), .C0(n31897), 
        .Y(n31899) );
  OAI211XL U34942 ( .A0(n35726), .A1(n31900), .B0(n16649), .C0(n31899), .Y(
        n15546) );
  NOR2BXL U34943 ( .AN(n31902), .B(n31901), .Y(n31904) );
  NAND2XL U34944 ( .A(conv_3[320]), .B(n31904), .Y(n31903) );
  OAI211XL U34945 ( .A0(conv_3[320]), .A1(n31904), .B0(n16656), .C0(n31903), 
        .Y(n31905) );
  OAI211XL U34946 ( .A0(n35743), .A1(n31906), .B0(n16649), .C0(n31905), .Y(
        n15533) );
  INVXL U34947 ( .A(conv_3[325]), .Y(n31914) );
  NOR2X1 U34948 ( .A(n33840), .B(n33281), .Y(n35739) );
  AOI21XL U34949 ( .A0(n31915), .A1(n33842), .B0(n31910), .Y(n31912) );
  NAND2XL U34950 ( .A(conv_3[325]), .B(n31912), .Y(n31911) );
  OAI211XL U34951 ( .A0(conv_3[325]), .A1(n31912), .B0(n32660), .C0(n31911), 
        .Y(n31913) );
  OAI211XL U34952 ( .A0(n35743), .A1(n31914), .B0(n33468), .C0(n31913), .Y(
        n15528) );
  OAI2BB1XL U34953 ( .A0N(conv_3[325]), .A1N(n31915), .B0(n33281), .Y(n33280)
         );
  NOR2X1 U34954 ( .A(conv_3[326]), .B(n31919), .Y(n33283) );
  AOI32XL U34955 ( .A0(conv_3[326]), .A1(n33281), .A2(n33280), .B0(n33842), 
        .B1(n33283), .Y(n31917) );
  NAND2XL U34956 ( .A(n33282), .B(n31917), .Y(n31916) );
  OAI211XL U34957 ( .A0(n33282), .A1(n31917), .B0(n33788), .C0(n31916), .Y(
        n31918) );
  OAI211XL U34958 ( .A0(n35743), .A1(n33282), .B0(n16649), .C0(n31918), .Y(
        n15526) );
  INVXL U34959 ( .A(conv_3[326]), .Y(n31923) );
  NAND2XL U34960 ( .A(conv_3[326]), .B(n31921), .Y(n31920) );
  OAI211XL U34961 ( .A0(conv_3[326]), .A1(n31921), .B0(n33822), .C0(n31920), 
        .Y(n31922) );
  OAI211XL U34962 ( .A0(n35743), .A1(n31923), .B0(n33468), .C0(n31922), .Y(
        n15527) );
  NAND2XL U34963 ( .A(conv_3[440]), .B(n31929), .Y(n31928) );
  OAI211XL U34964 ( .A0(conv_3[440]), .A1(n31929), .B0(n33788), .C0(n31928), 
        .Y(n31930) );
  OAI211XL U34965 ( .A0(n35792), .A1(n31931), .B0(n16649), .C0(n31930), .Y(
        n15453) );
  INVXL U34966 ( .A(conv_3[441]), .Y(n31937) );
  AOI2BB1XL U34967 ( .A0N(n33761), .A1N(n31939), .B0(n31938), .Y(n31935) );
  NAND2XL U34968 ( .A(conv_3[441]), .B(n31935), .Y(n31934) );
  OAI211XL U34969 ( .A0(conv_3[441]), .A1(n31935), .B0(n33788), .C0(n31934), 
        .Y(n31936) );
  OAI211XL U34970 ( .A0(n35792), .A1(n31937), .B0(n16649), .C0(n31936), .Y(
        n15452) );
  INVXL U34971 ( .A(conv_3[447]), .Y(n31944) );
  INVXL U34972 ( .A(conv_3[442]), .Y(n35784) );
  NAND2XL U34973 ( .A(conv_3[441]), .B(n31939), .Y(n35782) );
  NAND2XL U34974 ( .A(conv_3[443]), .B(n32110), .Y(n35788) );
  AOI21XL U34975 ( .A0(conv_3[445]), .A1(n33760), .B0(n33761), .Y(n31949) );
  AOI22XL U34976 ( .A0(n33761), .A1(n31945), .B0(n31943), .B1(n35789), .Y(
        n31941) );
  NAND2XL U34977 ( .A(n31944), .B(n31941), .Y(n31940) );
  OAI211XL U34978 ( .A0(n31944), .A1(n31941), .B0(n33778), .C0(n31940), .Y(
        n31942) );
  OAI211XL U34979 ( .A0(n35792), .A1(n31944), .B0(n16649), .C0(n31942), .Y(
        n15446) );
  NAND3XL U34980 ( .A(n31943), .B(conv_3[447]), .C(n35789), .Y(n32145) );
  NAND3XL U34981 ( .A(n31945), .B(n33761), .C(n31944), .Y(n32144) );
  NAND2XL U34982 ( .A(n32145), .B(n32144), .Y(n31947) );
  NAND2XL U34983 ( .A(conv_3[448]), .B(n31947), .Y(n31946) );
  OAI211XL U34984 ( .A0(conv_3[448]), .A1(n31947), .B0(n32611), .C0(n31946), 
        .Y(n31948) );
  OAI211XL U34985 ( .A0(n35792), .A1(n32143), .B0(n16649), .C0(n31948), .Y(
        n15445) );
  INVXL U34986 ( .A(conv_3[446]), .Y(n31954) );
  NAND2XL U34987 ( .A(conv_3[446]), .B(n31952), .Y(n31951) );
  OAI211XL U34988 ( .A0(conv_3[446]), .A1(n31952), .B0(n24378), .C0(n31951), 
        .Y(n31953) );
  OAI211XL U34989 ( .A0(n35792), .A1(n31954), .B0(n16649), .C0(n31953), .Y(
        n15447) );
  OAI21XL U34990 ( .A0(conv_3[340]), .A1(n31974), .B0(n31980), .Y(n31968) );
  NAND2XL U34991 ( .A(n31968), .B(n31981), .Y(n31959) );
  NAND2XL U34992 ( .A(n31969), .B(n31959), .Y(n31958) );
  OAI211XL U34993 ( .A0(n31969), .A1(n31959), .B0(n32660), .C0(n31958), .Y(
        n31960) );
  OAI211XL U34994 ( .A0(n35748), .A1(n31969), .B0(n16649), .C0(n31960), .Y(
        n15517) );
  INVXL U34995 ( .A(conv_3[338]), .Y(n31966) );
  AOI21XL U34996 ( .A0(n31962), .A1(n31980), .B0(n31961), .Y(n31964) );
  NAND2XL U34997 ( .A(conv_3[338]), .B(n31964), .Y(n31963) );
  OAI211XL U34998 ( .A0(conv_3[338]), .A1(n31964), .B0(n33712), .C0(n31963), 
        .Y(n31965) );
  OAI211XL U34999 ( .A0(n35748), .A1(n31966), .B0(n33468), .C0(n31965), .Y(
        n15520) );
  NAND4XL U35000 ( .A(conv_3[341]), .B(conv_3[342]), .C(n31967), .D(n31981), 
        .Y(n32215) );
  NAND2XL U35001 ( .A(n31969), .B(n31968), .Y(n31970) );
  NAND3XL U35002 ( .A(n31980), .B(n31986), .C(n31982), .Y(n32214) );
  NAND2XL U35003 ( .A(n32215), .B(n32214), .Y(n31972) );
  NAND2XL U35004 ( .A(conv_3[343]), .B(n31972), .Y(n31971) );
  OAI211XL U35005 ( .A0(conv_3[343]), .A1(n31972), .B0(n36020), .C0(n31971), 
        .Y(n31973) );
  OAI211XL U35006 ( .A0(n35748), .A1(n32213), .B0(n16649), .C0(n31973), .Y(
        n15515) );
  INVXL U35007 ( .A(conv_3[340]), .Y(n31979) );
  NAND2XL U35008 ( .A(conv_3[340]), .B(n31977), .Y(n31976) );
  OAI211XL U35009 ( .A0(conv_3[340]), .A1(n31977), .B0(n33982), .C0(n31976), 
        .Y(n31978) );
  OAI211XL U35010 ( .A0(n35748), .A1(n31979), .B0(n33468), .C0(n31978), .Y(
        n15518) );
  AOI32XL U35011 ( .A0(conv_3[341]), .A1(n31982), .A2(n31981), .B0(n31980), 
        .B1(n31982), .Y(n31984) );
  NAND2XL U35012 ( .A(n31986), .B(n31984), .Y(n31983) );
  OAI211XL U35013 ( .A0(n31986), .A1(n31984), .B0(n31735), .C0(n31983), .Y(
        n31985) );
  OAI211XL U35014 ( .A0(n35748), .A1(n31986), .B0(n16649), .C0(n31985), .Y(
        n15516) );
  NOR2BXL U35015 ( .AN(n31988), .B(n31987), .Y(n31990) );
  NAND2XL U35016 ( .A(conv_3[412]), .B(n31990), .Y(n31989) );
  OAI211XL U35017 ( .A0(conv_3[412]), .A1(n31990), .B0(n33822), .C0(n31989), 
        .Y(n31991) );
  OAI211XL U35018 ( .A0(n34227), .A1(n31992), .B0(n16649), .C0(n31991), .Y(
        n15471) );
  INVXL U35019 ( .A(conv_3[417]), .Y(n32000) );
  AOI31XL U35020 ( .A0(conv_3[415]), .A1(conv_3[414]), .A2(n32559), .B0(n32557), .Y(n32010) );
  OAI21XL U35021 ( .A0(n32557), .A1(n31998), .B0(n31999), .Y(n31996) );
  NAND2XL U35022 ( .A(n32000), .B(n31996), .Y(n31995) );
  OAI211XL U35023 ( .A0(n32000), .A1(n31996), .B0(n24499), .C0(n31995), .Y(
        n31997) );
  OAI211XL U35024 ( .A0(n34227), .A1(n32000), .B0(n33468), .C0(n31997), .Y(
        n15466) );
  NAND3XL U35025 ( .A(n31998), .B(conv_3[417]), .C(n32558), .Y(n32192) );
  NAND3XL U35026 ( .A(n32557), .B(n32000), .C(n31999), .Y(n32191) );
  NAND2XL U35027 ( .A(n32192), .B(n32191), .Y(n32002) );
  NAND2XL U35028 ( .A(conv_3[418]), .B(n32002), .Y(n32001) );
  OAI211XL U35029 ( .A0(conv_3[418]), .A1(n32002), .B0(n33788), .C0(n32001), 
        .Y(n32003) );
  OAI211XL U35030 ( .A0(n34227), .A1(n32190), .B0(n16649), .C0(n32003), .Y(
        n15465) );
  INVXL U35031 ( .A(conv_3[411]), .Y(n32009) );
  AOI2BB1XL U35032 ( .A0N(n32557), .A1N(n32005), .B0(n32004), .Y(n32007) );
  NAND2XL U35033 ( .A(conv_3[411]), .B(n32007), .Y(n32006) );
  OAI211XL U35034 ( .A0(conv_3[411]), .A1(n32007), .B0(n33788), .C0(n32006), 
        .Y(n32008) );
  OAI211XL U35035 ( .A0(n34227), .A1(n32009), .B0(n33468), .C0(n32008), .Y(
        n15472) );
  NAND2XL U35036 ( .A(conv_3[416]), .B(n32013), .Y(n32012) );
  OAI211XL U35037 ( .A0(conv_3[416]), .A1(n32013), .B0(n16657), .C0(n32012), 
        .Y(n32014) );
  OAI211XL U35038 ( .A0(n34227), .A1(n32015), .B0(n33468), .C0(n32014), .Y(
        n15467) );
  INVXL U35039 ( .A(conv_3[395]), .Y(n32024) );
  NAND2XL U35040 ( .A(conv_3[395]), .B(n32022), .Y(n32021) );
  OAI211XL U35041 ( .A0(conv_3[395]), .A1(n32022), .B0(n32052), .C0(n32021), 
        .Y(n32023) );
  OAI211XL U35042 ( .A0(n33703), .A1(n32024), .B0(n16649), .C0(n32023), .Y(
        n15483) );
  INVXL U35043 ( .A(conv_3[396]), .Y(n32030) );
  INVXL U35044 ( .A(n33699), .Y(n33695) );
  AOI2BB1XL U35045 ( .A0N(n33699), .A1N(n32031), .B0(n32032), .Y(n32028) );
  NAND2XL U35046 ( .A(conv_3[396]), .B(n32028), .Y(n32027) );
  OAI211XL U35047 ( .A0(conv_3[396]), .A1(n32028), .B0(n32052), .C0(n32027), 
        .Y(n32029) );
  OAI211XL U35048 ( .A0(n33703), .A1(n32030), .B0(n16649), .C0(n32029), .Y(
        n15482) );
  INVXL U35049 ( .A(conv_3[397]), .Y(n32036) );
  AOI21XL U35050 ( .A0(n32031), .A1(conv_3[396]), .B0(n33699), .Y(n32037) );
  NAND2XL U35051 ( .A(conv_3[397]), .B(n32034), .Y(n32033) );
  OAI211XL U35052 ( .A0(conv_3[397]), .A1(n32034), .B0(n32052), .C0(n32033), 
        .Y(n32035) );
  OAI211XL U35053 ( .A0(n33703), .A1(n32036), .B0(n33468), .C0(n32035), .Y(
        n15481) );
  NAND2XL U35054 ( .A(n33699), .B(n32048), .Y(n32043) );
  NAND2XL U35055 ( .A(n32047), .B(n32043), .Y(n32050) );
  AOI31XL U35056 ( .A0(conv_3[400]), .A1(conv_3[399]), .A2(n32048), .B0(n33699), .Y(n33221) );
  NAND2XL U35057 ( .A(conv_3[401]), .B(n32040), .Y(n32039) );
  OAI211XL U35058 ( .A0(conv_3[401]), .A1(n32040), .B0(n33982), .C0(n32039), 
        .Y(n32041) );
  OAI211XL U35059 ( .A0(n33703), .A1(n32042), .B0(n33468), .C0(n32041), .Y(
        n15477) );
  OAI21XL U35060 ( .A0(n33699), .A1(n32048), .B0(n32043), .Y(n32045) );
  NAND2XL U35061 ( .A(n32047), .B(n32045), .Y(n32044) );
  OAI211XL U35062 ( .A0(n32047), .A1(n32045), .B0(n32052), .C0(n32044), .Y(
        n32046) );
  OAI211XL U35063 ( .A0(n33703), .A1(n32047), .B0(n33468), .C0(n32046), .Y(
        n15479) );
  INVXL U35064 ( .A(conv_3[400]), .Y(n32055) );
  AOI21XL U35065 ( .A0(conv_3[399]), .A1(n32048), .B0(n33699), .Y(n32049) );
  AOI21XL U35066 ( .A0(n33699), .A1(n32050), .B0(n32049), .Y(n32053) );
  NAND2XL U35067 ( .A(conv_3[400]), .B(n32053), .Y(n32051) );
  OAI211XL U35068 ( .A0(conv_3[400]), .A1(n32053), .B0(n32052), .C0(n32051), 
        .Y(n32054) );
  OAI211XL U35069 ( .A0(n33703), .A1(n32055), .B0(n33468), .C0(n32054), .Y(
        n15478) );
  AOI221XL U35070 ( .A0(n32057), .A1(n33778), .B0(n32056), .B1(n16657), .C0(
        n35662), .Y(n32062) );
  OAI211XL U35071 ( .A0(n35660), .A1(n32059), .B0(n33912), .C0(n32058), .Y(
        n32060) );
  OAI211XL U35072 ( .A0(n32062), .A1(n32061), .B0(n33468), .C0(n32060), .Y(
        n15600) );
  INVXL U35073 ( .A(conv_3[505]), .Y(n32069) );
  NAND2XL U35074 ( .A(conv_3[503]), .B(n32083), .Y(n32077) );
  AOI2BB1XL U35075 ( .A0N(n35838), .A1N(n32346), .B0(n32345), .Y(n32067) );
  NAND2XL U35076 ( .A(conv_3[505]), .B(n32067), .Y(n32066) );
  OAI211XL U35077 ( .A0(conv_3[505]), .A1(n32067), .B0(n33788), .C0(n32066), 
        .Y(n32068) );
  OAI211XL U35078 ( .A0(n35841), .A1(n32069), .B0(n16649), .C0(n32068), .Y(
        n15408) );
  NAND2XL U35079 ( .A(conv_3[500]), .B(n32073), .Y(n32072) );
  OAI211XL U35080 ( .A0(conv_3[500]), .A1(n32073), .B0(n33982), .C0(n32072), 
        .Y(n32074) );
  OAI211XL U35081 ( .A0(n35841), .A1(n32075), .B0(n16649), .C0(n32074), .Y(
        n15413) );
  AOI21XL U35082 ( .A0(n33918), .A1(n32077), .B0(n32076), .Y(n32079) );
  NAND2XL U35083 ( .A(conv_3[504]), .B(n32079), .Y(n32078) );
  OAI211XL U35084 ( .A0(conv_3[504]), .A1(n32079), .B0(n31735), .C0(n32078), 
        .Y(n32080) );
  OAI211XL U35085 ( .A0(n35841), .A1(n32081), .B0(n16649), .C0(n32080), .Y(
        n15409) );
  INVXL U35086 ( .A(conv_3[503]), .Y(n32087) );
  AOI2BB1XL U35087 ( .A0N(n35838), .A1N(n32083), .B0(n32082), .Y(n32085) );
  NAND2XL U35088 ( .A(conv_3[503]), .B(n32085), .Y(n32084) );
  OAI211XL U35089 ( .A0(conv_3[503]), .A1(n32085), .B0(n27932), .C0(n32084), 
        .Y(n32086) );
  OAI211XL U35090 ( .A0(n35841), .A1(n32087), .B0(n16649), .C0(n32086), .Y(
        n15410) );
  AOI2BB1XL U35091 ( .A0N(n35673), .A1N(n32089), .B0(n32088), .Y(n32091) );
  NAND2XL U35092 ( .A(conv_3[231]), .B(n32091), .Y(n32090) );
  OAI211XL U35093 ( .A0(conv_3[231]), .A1(n32091), .B0(n33912), .C0(n32090), 
        .Y(n32092) );
  OAI211XL U35094 ( .A0(n35676), .A1(n32093), .B0(n33468), .C0(n32092), .Y(
        n15592) );
  AOI21XL U35095 ( .A0(n33878), .A1(n32095), .B0(n32094), .Y(n32097) );
  NAND2XL U35096 ( .A(conv_3[232]), .B(n32097), .Y(n32096) );
  OAI211XL U35097 ( .A0(conv_3[232]), .A1(n32097), .B0(n33912), .C0(n32096), 
        .Y(n32098) );
  OAI211XL U35098 ( .A0(n35676), .A1(n32099), .B0(n33468), .C0(n32098), .Y(
        n15591) );
  AOI2BB1XL U35099 ( .A0N(n33480), .A1N(n33006), .B0(n33007), .Y(n32104) );
  NAND2XL U35100 ( .A(conv_3[264]), .B(n32104), .Y(n32103) );
  OAI211XL U35101 ( .A0(conv_3[264]), .A1(n32104), .B0(n31735), .C0(n32103), 
        .Y(n32105) );
  OAI211XL U35102 ( .A0(n35713), .A1(n32106), .B0(n16649), .C0(n32105), .Y(
        n15569) );
  AOI221XL U35103 ( .A0(n32108), .A1(n32052), .B0(n32107), .B1(n35336), .C0(
        n33756), .Y(n32113) );
  OAI211XL U35104 ( .A0(n33761), .A1(n32110), .B0(n16657), .C0(n32109), .Y(
        n32111) );
  OAI211XL U35105 ( .A0(n32113), .A1(n32112), .B0(n16649), .C0(n32111), .Y(
        n15450) );
  OAI2BB1XL U35106 ( .A0N(conv_3[100]), .A1N(n32114), .B0(n35615), .Y(n34187)
         );
  NAND4XL U35107 ( .A(conv_3[101]), .B(conv_3[102]), .C(n35615), .D(n34187), 
        .Y(n32666) );
  INVXL U35108 ( .A(conv_3[101]), .Y(n34184) );
  OAI21XL U35109 ( .A0(conv_3[100]), .A1(n32115), .B0(n34186), .Y(n34180) );
  NAND2XL U35110 ( .A(n34184), .B(n34180), .Y(n32116) );
  NAND3XL U35111 ( .A(n34186), .B(n34192), .C(n34188), .Y(n32665) );
  INVXL U35112 ( .A(conv_3[103]), .Y(n32669) );
  AOI22XL U35113 ( .A0(conv_3[103]), .A1(n32666), .B0(n32665), .B1(n32669), 
        .Y(n32118) );
  NAND2XL U35114 ( .A(conv_3[104]), .B(n32118), .Y(n32117) );
  OAI211XL U35115 ( .A0(conv_3[104]), .A1(n32118), .B0(n32052), .C0(n32117), 
        .Y(n32119) );
  OAI211XL U35116 ( .A0(n34789), .A1(n32120), .B0(n33468), .C0(n32119), .Y(
        n15674) );
  AOI22XL U35117 ( .A0(conv_3[373]), .A1(n32123), .B0(n32122), .B1(n32121), 
        .Y(n32125) );
  NAND2XL U35118 ( .A(conv_3[374]), .B(n32125), .Y(n32124) );
  OAI211XL U35119 ( .A0(conv_3[374]), .A1(n32125), .B0(n16657), .C0(n32124), 
        .Y(n32126) );
  OAI211XL U35120 ( .A0(n34520), .A1(n32127), .B0(n33468), .C0(n32126), .Y(
        n15494) );
  NAND3XL U35121 ( .A(n33726), .B(conv_3[357]), .C(n32130), .Y(n34745) );
  NAND2XL U35122 ( .A(n33752), .B(n33725), .Y(n34744) );
  AOI22XL U35123 ( .A0(conv_3[358]), .A1(n34745), .B0(n34744), .B1(n34749), 
        .Y(n32133) );
  NAND2XL U35124 ( .A(conv_3[359]), .B(n32133), .Y(n32132) );
  OAI211XL U35125 ( .A0(conv_3[359]), .A1(n32133), .B0(n24378), .C0(n32132), 
        .Y(n32134) );
  OAI211XL U35126 ( .A0(n34520), .A1(n32135), .B0(n16649), .C0(n32134), .Y(
        n15504) );
  AOI22XL U35127 ( .A0(conv_3[223]), .A1(n32138), .B0(n32137), .B1(n32136), 
        .Y(n32140) );
  NAND2XL U35128 ( .A(conv_3[224]), .B(n32140), .Y(n32139) );
  OAI211XL U35129 ( .A0(conv_3[224]), .A1(n32140), .B0(n33912), .C0(n32139), 
        .Y(n32141) );
  OAI211XL U35130 ( .A0(n34520), .A1(n32142), .B0(n33468), .C0(n32141), .Y(
        n15594) );
  AOI22XL U35131 ( .A0(conv_3[448]), .A1(n32145), .B0(n32144), .B1(n32143), 
        .Y(n32147) );
  NAND2XL U35132 ( .A(conv_3[449]), .B(n32147), .Y(n32146) );
  OAI211XL U35133 ( .A0(conv_3[449]), .A1(n32147), .B0(n35336), .C0(n32146), 
        .Y(n32148) );
  OAI211XL U35134 ( .A0(n34520), .A1(n32149), .B0(n16649), .C0(n32148), .Y(
        n15444) );
  AOI22XL U35135 ( .A0(conv_3[88]), .A1(n32152), .B0(n32151), .B1(n32150), .Y(
        n32154) );
  NAND2XL U35136 ( .A(conv_3[89]), .B(n32154), .Y(n32153) );
  OAI211XL U35137 ( .A0(conv_3[89]), .A1(n32154), .B0(n33788), .C0(n32153), 
        .Y(n32155) );
  OAI211XL U35138 ( .A0(n34789), .A1(n32156), .B0(n33468), .C0(n32155), .Y(
        n15684) );
  NAND4XL U35139 ( .A(conv_3[431]), .B(conv_3[432]), .C(n35775), .D(n32582), 
        .Y(n32588) );
  INVXL U35140 ( .A(n32581), .Y(n32158) );
  AOI21XL U35141 ( .A0(conv_3[433]), .A1(n32588), .B0(n32589), .Y(n32160) );
  NAND2XL U35142 ( .A(conv_3[434]), .B(n32160), .Y(n32159) );
  OAI211XL U35143 ( .A0(conv_3[434]), .A1(n32160), .B0(n34028), .C0(n32159), 
        .Y(n32161) );
  OAI211XL U35144 ( .A0(n34520), .A1(n32162), .B0(n16649), .C0(n32161), .Y(
        n15454) );
  NAND3XL U35145 ( .A(conv_3[72]), .B(n32164), .C(n32163), .Y(n32570) );
  OR3XL U35146 ( .A(n32164), .B(conv_3[72]), .C(n32163), .Y(n32569) );
  INVXL U35147 ( .A(conv_3[73]), .Y(n32573) );
  AOI22XL U35148 ( .A0(conv_3[73]), .A1(n32570), .B0(n32569), .B1(n32573), .Y(
        n32166) );
  NAND2XL U35149 ( .A(conv_3[74]), .B(n32166), .Y(n32165) );
  OAI211XL U35150 ( .A0(conv_3[74]), .A1(n32166), .B0(n33778), .C0(n32165), 
        .Y(n32167) );
  AOI22XL U35151 ( .A0(conv_3[148]), .A1(n32171), .B0(n32170), .B1(n32169), 
        .Y(n32173) );
  NAND2XL U35152 ( .A(conv_3[149]), .B(n32173), .Y(n32172) );
  OAI211XL U35153 ( .A0(conv_3[149]), .A1(n32173), .B0(n36020), .C0(n32172), 
        .Y(n32174) );
  OAI211XL U35154 ( .A0(n34789), .A1(n32175), .B0(n33468), .C0(n32174), .Y(
        n15644) );
  NAND3XL U35155 ( .A(n33823), .B(conv_3[57]), .C(n32178), .Y(n34157) );
  NAND2XL U35156 ( .A(n33824), .B(n33821), .Y(n34156) );
  AOI22XL U35157 ( .A0(conv_3[58]), .A1(n34157), .B0(n34156), .B1(n34160), .Y(
        n32182) );
  NAND2XL U35158 ( .A(conv_3[59]), .B(n32182), .Y(n32180) );
  OAI211XL U35159 ( .A0(conv_3[59]), .A1(n32182), .B0(n32181), .C0(n32180), 
        .Y(n32183) );
  OAI211XL U35160 ( .A0(n34789), .A1(n32184), .B0(n33468), .C0(n32183), .Y(
        n15704) );
  NAND4XL U35161 ( .A(conv_3[476]), .B(conv_3[477]), .C(n32328), .D(n32340), 
        .Y(n32322) );
  NAND3XL U35162 ( .A(n32327), .B(n35810), .C(n32332), .Y(n32321) );
  OAI211XL U35163 ( .A0(conv_3[479]), .A1(n32187), .B0(n34028), .C0(n32186), 
        .Y(n32188) );
  OAI211XL U35164 ( .A0(n34520), .A1(n32189), .B0(n16649), .C0(n32188), .Y(
        n15424) );
  AOI22XL U35165 ( .A0(conv_3[418]), .A1(n32192), .B0(n32191), .B1(n32190), 
        .Y(n32194) );
  NAND2XL U35166 ( .A(conv_3[419]), .B(n32194), .Y(n32193) );
  OAI211XL U35167 ( .A0(conv_3[419]), .A1(n32194), .B0(n24499), .C0(n32193), 
        .Y(n32195) );
  OAI211XL U35168 ( .A0(n34520), .A1(n32196), .B0(n16649), .C0(n32195), .Y(
        n15464) );
  NAND3XL U35169 ( .A(n34163), .B(conv_3[387]), .C(n32200), .Y(n34139) );
  AOI22XL U35170 ( .A0(conv_3[388]), .A1(n34139), .B0(n34138), .B1(n34142), 
        .Y(n32202) );
  NAND2XL U35171 ( .A(conv_3[389]), .B(n32202), .Y(n32201) );
  OAI211XL U35172 ( .A0(conv_3[389]), .A1(n32202), .B0(n33778), .C0(n32201), 
        .Y(n32203) );
  NAND2XL U35173 ( .A(conv_3[194]), .B(n32210), .Y(n32209) );
  OAI211XL U35174 ( .A0(conv_3[194]), .A1(n32210), .B0(n33912), .C0(n32209), 
        .Y(n32211) );
  OAI211XL U35175 ( .A0(n34676), .A1(n32212), .B0(n33468), .C0(n32211), .Y(
        n15614) );
  AOI22XL U35176 ( .A0(conv_3[343]), .A1(n32215), .B0(n32214), .B1(n32213), 
        .Y(n32217) );
  NAND2XL U35177 ( .A(conv_3[344]), .B(n32217), .Y(n32216) );
  OAI211XL U35178 ( .A0(conv_3[344]), .A1(n32217), .B0(n33712), .C0(n32216), 
        .Y(n32218) );
  OAI211XL U35179 ( .A0(n34789), .A1(n32219), .B0(n16649), .C0(n32218), .Y(
        n15514) );
  NAND3XL U35180 ( .A(conv_3[177]), .B(n32220), .C(n32221), .Y(n32642) );
  AOI21XL U35181 ( .A0(conv_3[178]), .A1(n32642), .B0(n32643), .Y(n32224) );
  NAND2XL U35182 ( .A(conv_3[179]), .B(n32224), .Y(n32223) );
  OAI211XL U35183 ( .A0(conv_3[179]), .A1(n32224), .B0(n34028), .C0(n32223), 
        .Y(n32225) );
  OAI211XL U35184 ( .A0(n34789), .A1(n32226), .B0(n33468), .C0(n32225), .Y(
        n15624) );
  NAND4XL U35185 ( .A(conv_3[491]), .B(conv_3[492]), .C(n35823), .D(n32227), 
        .Y(n33309) );
  NAND3XL U35186 ( .A(n35831), .B(n32229), .C(n32228), .Y(n33308) );
  INVXL U35187 ( .A(conv_3[493]), .Y(n33312) );
  AOI22XL U35188 ( .A0(conv_3[493]), .A1(n33309), .B0(n33308), .B1(n33312), 
        .Y(n32231) );
  NAND2XL U35189 ( .A(conv_3[494]), .B(n32231), .Y(n32230) );
  OAI211XL U35190 ( .A0(conv_3[494]), .A1(n32231), .B0(n31735), .C0(n32230), 
        .Y(n32232) );
  OAI211XL U35191 ( .A0(n34520), .A1(n32233), .B0(n16649), .C0(n32232), .Y(
        n15414) );
  AOI22XL U35192 ( .A0(conv_3[298]), .A1(n32236), .B0(n32235), .B1(n32234), 
        .Y(n32238) );
  NAND2XL U35193 ( .A(conv_3[299]), .B(n32238), .Y(n32237) );
  OAI211XL U35194 ( .A0(conv_3[299]), .A1(n32238), .B0(n34666), .C0(n32237), 
        .Y(n32239) );
  OAI211XL U35195 ( .A0(n34789), .A1(n32240), .B0(n16649), .C0(n32239), .Y(
        n15544) );
  AOI22XL U35196 ( .A0(conv_3[463]), .A1(n32243), .B0(n32242), .B1(n32241), 
        .Y(n32245) );
  NAND2XL U35197 ( .A(conv_3[464]), .B(n32245), .Y(n32244) );
  OAI211XL U35198 ( .A0(conv_3[464]), .A1(n32245), .B0(n33712), .C0(n32244), 
        .Y(n32246) );
  OAI211XL U35199 ( .A0(n34520), .A1(n32247), .B0(n16649), .C0(n32246), .Y(
        n15434) );
  AOI21XL U35200 ( .A0(conv_3[158]), .A1(n32279), .B0(n32316), .Y(n32296) );
  NAND3XL U35201 ( .A(n32291), .B(conv_3[162]), .C(n32252), .Y(n34468) );
  INVXL U35202 ( .A(conv_3[160]), .Y(n32307) );
  NAND2XL U35203 ( .A(n32307), .B(n32302), .Y(n32315) );
  OAI21XL U35204 ( .A0(conv_3[161]), .A1(n32315), .B0(n32316), .Y(n32290) );
  NAND3XL U35205 ( .A(n32316), .B(n32295), .C(n32290), .Y(n34467) );
  INVXL U35206 ( .A(conv_3[163]), .Y(n34471) );
  AOI22XL U35207 ( .A0(conv_3[163]), .A1(n34468), .B0(n34467), .B1(n34471), 
        .Y(n32254) );
  NAND2XL U35208 ( .A(conv_3[164]), .B(n32254), .Y(n32253) );
  OAI211XL U35209 ( .A0(conv_3[164]), .A1(n32254), .B0(n32052), .C0(n32253), 
        .Y(n32255) );
  OAI211XL U35210 ( .A0(n34789), .A1(n32256), .B0(n33468), .C0(n32255), .Y(
        n15634) );
  AOI22XL U35211 ( .A0(conv_3[283]), .A1(n32259), .B0(n32258), .B1(n32257), 
        .Y(n32261) );
  NAND2XL U35212 ( .A(conv_3[284]), .B(n32261), .Y(n32260) );
  OAI211XL U35213 ( .A0(conv_3[284]), .A1(n32261), .B0(n35336), .C0(n32260), 
        .Y(n32262) );
  OAI211XL U35214 ( .A0(n34789), .A1(n32263), .B0(n16649), .C0(n32262), .Y(
        n15554) );
  AOI22XL U35215 ( .A0(conv_3[118]), .A1(n32266), .B0(n32265), .B1(n32264), 
        .Y(n32268) );
  NAND2XL U35216 ( .A(conv_3[119]), .B(n32268), .Y(n32267) );
  OAI211XL U35217 ( .A0(conv_3[119]), .A1(n32268), .B0(n34028), .C0(n32267), 
        .Y(n32269) );
  OAI211XL U35218 ( .A0(n34789), .A1(n32270), .B0(n16649), .C0(n32269), .Y(
        n15664) );
  AOI22XL U35219 ( .A0(conv_3[208]), .A1(n32273), .B0(n32272), .B1(n32271), 
        .Y(n32275) );
  NAND2XL U35220 ( .A(conv_3[209]), .B(n32275), .Y(n32274) );
  OAI211XL U35221 ( .A0(conv_3[209]), .A1(n32275), .B0(n33912), .C0(n32274), 
        .Y(n32276) );
  OAI211XL U35222 ( .A0(n34520), .A1(n32277), .B0(n33468), .C0(n32276), .Y(
        n15604) );
  INVXL U35223 ( .A(conv_3[158]), .Y(n32283) );
  AOI2BB1XL U35224 ( .A0N(n32316), .A1N(n32279), .B0(n32278), .Y(n32281) );
  NAND2XL U35225 ( .A(conv_3[158]), .B(n32281), .Y(n32280) );
  OAI211XL U35226 ( .A0(conv_3[158]), .A1(n32281), .B0(n34666), .C0(n32280), 
        .Y(n32282) );
  OAI211XL U35227 ( .A0(n34751), .A1(n32283), .B0(n33468), .C0(n32282), .Y(
        n15640) );
  NAND2XL U35228 ( .A(conv_3[155]), .B(n32287), .Y(n32286) );
  OAI211XL U35229 ( .A0(conv_3[155]), .A1(n32287), .B0(n31735), .C0(n32286), 
        .Y(n32288) );
  OAI211XL U35230 ( .A0(n34751), .A1(n32289), .B0(n33468), .C0(n32288), .Y(
        n15643) );
  OAI21XL U35231 ( .A0(n32316), .A1(n32291), .B0(n32290), .Y(n32293) );
  NAND2XL U35232 ( .A(n32295), .B(n32293), .Y(n32292) );
  OAI211XL U35233 ( .A0(n32295), .A1(n32293), .B0(n32052), .C0(n32292), .Y(
        n32294) );
  OAI211XL U35234 ( .A0(n34751), .A1(n32295), .B0(n33468), .C0(n32294), .Y(
        n15636) );
  INVXL U35235 ( .A(conv_3[159]), .Y(n32301) );
  NAND2XL U35236 ( .A(conv_3[159]), .B(n32299), .Y(n32298) );
  OAI211XL U35237 ( .A0(conv_3[159]), .A1(n32299), .B0(n33778), .C0(n32298), 
        .Y(n32300) );
  OAI211XL U35238 ( .A0(n34751), .A1(n32301), .B0(n33468), .C0(n32300), .Y(
        n15639) );
  OAI21XL U35239 ( .A0(n32316), .A1(n32303), .B0(n32302), .Y(n32305) );
  NAND2XL U35240 ( .A(n32307), .B(n32305), .Y(n32304) );
  OAI211XL U35241 ( .A0(n32307), .A1(n32305), .B0(n33778), .C0(n32304), .Y(
        n32306) );
  OAI211XL U35242 ( .A0(n34751), .A1(n32307), .B0(n33468), .C0(n32306), .Y(
        n15638) );
  AOI2BB1XL U35243 ( .A0N(n32316), .A1N(n32309), .B0(n32308), .Y(n32311) );
  NAND2XL U35244 ( .A(conv_3[156]), .B(n32311), .Y(n32310) );
  OAI211XL U35245 ( .A0(conv_3[156]), .A1(n32311), .B0(n28751), .C0(n32310), 
        .Y(n32312) );
  OAI211XL U35246 ( .A0(n34751), .A1(n32313), .B0(n33468), .C0(n32312), .Y(
        n15642) );
  AOI21XL U35247 ( .A0(n32316), .A1(n32315), .B0(n32314), .Y(n32318) );
  NAND2XL U35248 ( .A(conv_3[161]), .B(n32318), .Y(n32317) );
  OAI211XL U35249 ( .A0(conv_3[161]), .A1(n32318), .B0(n33788), .C0(n32317), 
        .Y(n32319) );
  OAI211XL U35250 ( .A0(n34751), .A1(n32320), .B0(n33468), .C0(n32319), .Y(
        n15637) );
  NAND2XL U35251 ( .A(n32322), .B(n32321), .Y(n32324) );
  NAND2XL U35252 ( .A(conv_3[478]), .B(n32324), .Y(n32323) );
  OAI211XL U35253 ( .A0(conv_3[478]), .A1(n32324), .B0(n32611), .C0(n32323), 
        .Y(n32325) );
  OAI211XL U35254 ( .A0(n35813), .A1(n32326), .B0(n16649), .C0(n32325), .Y(
        n15425) );
  AOI32XL U35255 ( .A0(conv_3[476]), .A1(n32328), .A2(n32340), .B0(n35810), 
        .B1(n32327), .Y(n32330) );
  NAND2XL U35256 ( .A(n32332), .B(n32330), .Y(n32329) );
  OAI211XL U35257 ( .A0(n32332), .A1(n32330), .B0(n32181), .C0(n32329), .Y(
        n32331) );
  OAI211XL U35258 ( .A0(n35813), .A1(n32332), .B0(n16649), .C0(n32331), .Y(
        n15426) );
  NAND2XL U35259 ( .A(conv_3[472]), .B(n32336), .Y(n32335) );
  OAI211XL U35260 ( .A0(conv_3[472]), .A1(n32336), .B0(n33157), .C0(n32335), 
        .Y(n32337) );
  OAI211XL U35261 ( .A0(n35813), .A1(n32338), .B0(n16649), .C0(n32337), .Y(
        n15431) );
  NAND2XL U35262 ( .A(conv_3[476]), .B(n32342), .Y(n32341) );
  OAI211XL U35263 ( .A0(conv_3[476]), .A1(n32342), .B0(n16656), .C0(n32341), 
        .Y(n32343) );
  OAI211XL U35264 ( .A0(n35813), .A1(n32344), .B0(n16649), .C0(n32343), .Y(
        n15427) );
  INVXL U35265 ( .A(conv_3[506]), .Y(n33855) );
  OAI21XL U35266 ( .A0(conv_3[505]), .A1(n32345), .B0(n35838), .Y(n33854) );
  OAI2BB1XL U35267 ( .A0N(conv_3[505]), .A1N(n32346), .B0(n33918), .Y(n33917)
         );
  NAND2XL U35268 ( .A(n33854), .B(n33917), .Y(n32348) );
  NAND2XL U35269 ( .A(n33855), .B(n32348), .Y(n32347) );
  OAI211XL U35270 ( .A0(n33855), .A1(n32348), .B0(n33788), .C0(n32347), .Y(
        n32349) );
  OAI211XL U35271 ( .A0(n35841), .A1(n33855), .B0(n16649), .C0(n32349), .Y(
        n15407) );
  INVXL U35272 ( .A(weight_1[25]), .Y(n32352) );
  OAI22XL U35273 ( .A0(n16650), .A1(n32352), .B0(n32350), .B1(n26910), .Y(
        n14434) );
  INVXL U35274 ( .A(weight_1[115]), .Y(n32353) );
  INVXL U35275 ( .A(weight_1[121]), .Y(n32357) );
  OAI22XL U35276 ( .A0(n16650), .A1(n32353), .B0(n32357), .B1(n26910), .Y(
        n14449) );
  INVXL U35277 ( .A(weight_1[7]), .Y(n32364) );
  OAI22XL U35278 ( .A0(n26906), .A1(n32351), .B0(n32364), .B1(n26910), .Y(
        n14430) );
  INVXL U35279 ( .A(weight_1[19]), .Y(n32359) );
  OAI22XL U35280 ( .A0(n31071), .A1(n32359), .B0(n32352), .B1(n26910), .Y(
        n14433) );
  OAI22XL U35281 ( .A0(n31077), .A1(n32354), .B0(n32353), .B1(n26910), .Y(
        n14448) );
  INVXL U35282 ( .A(weight_1[464]), .Y(n32358) );
  OAI22XL U35283 ( .A0(n31077), .A1(n32358), .B0(n32355), .B1(n16647), .Y(
        n14426) );
  INVXL U35284 ( .A(weight_1[97]), .Y(n32360) );
  OAI22XL U35285 ( .A0(n31084), .A1(n32360), .B0(n32356), .B1(n26910), .Y(
        n14446) );
  INVXL U35286 ( .A(weight_1[127]), .Y(n32482) );
  OAI22XL U35287 ( .A0(n32491), .A1(n32357), .B0(n32482), .B1(n16647), .Y(
        n14450) );
  OAI22XL U35288 ( .A0(n16650), .A1(n32372), .B0(n32358), .B1(n26910), .Y(
        n14425) );
  INVXL U35289 ( .A(weight_1[79]), .Y(n32685) );
  INVXL U35290 ( .A(weight_1[85]), .Y(n32362) );
  OAI22XL U35291 ( .A0(n31077), .A1(n32685), .B0(n32362), .B1(n26910), .Y(
        n14443) );
  INVXL U35292 ( .A(weight_1[13]), .Y(n32363) );
  OAI22XL U35293 ( .A0(n32967), .A1(n32363), .B0(n32359), .B1(n26910), .Y(
        n14432) );
  INVXL U35294 ( .A(weight_1[91]), .Y(n32361) );
  OAI22XL U35295 ( .A0(n31077), .A1(n32361), .B0(n32360), .B1(n16646), .Y(
        n14445) );
  OAI22XL U35296 ( .A0(n16650), .A1(n32362), .B0(n32361), .B1(n26910), .Y(
        n14444) );
  INVXL U35297 ( .A(weight_1[49]), .Y(n32680) );
  INVXL U35298 ( .A(weight_1[55]), .Y(n32682) );
  OAI22XL U35299 ( .A0(n16650), .A1(n32680), .B0(n32682), .B1(n26910), .Y(
        n14438) );
  OAI22XL U35300 ( .A0(n32491), .A1(n32364), .B0(n32363), .B1(n26910), .Y(
        n14431) );
  OAI22XL U35301 ( .A0(n16650), .A1(n32678), .B0(n36142), .B1(n16647), .Y(
        n14429) );
  INVXL U35302 ( .A(weight_1[308]), .Y(n32712) );
  INVXL U35303 ( .A(weight_1[314]), .Y(n32722) );
  OAI22XL U35304 ( .A0(n32491), .A1(n32712), .B0(n32722), .B1(n16646), .Y(
        n14400) );
  INVXL U35305 ( .A(weight_1[14]), .Y(n32377) );
  OAI22XL U35306 ( .A0(n32491), .A1(n32377), .B0(n32365), .B1(n16647), .Y(
        n14351) );
  INVXL U35307 ( .A(weight_1[362]), .Y(n32716) );
  INVXL U35308 ( .A(weight_1[368]), .Y(n32374) );
  OAI22XL U35309 ( .A0(n32491), .A1(n32716), .B0(n32374), .B1(n16646), .Y(
        n14409) );
  INVXL U35310 ( .A(weight_1[110]), .Y(n32393) );
  INVXL U35311 ( .A(weight_1[116]), .Y(n32708) );
  OAI22XL U35312 ( .A0(n16645), .A1(n32393), .B0(n32708), .B1(n16647), .Y(
        n14367) );
  INVXL U35313 ( .A(weight_1[416]), .Y(n32395) );
  OAI22XL U35314 ( .A0(n31077), .A1(n32395), .B0(n32366), .B1(n16646), .Y(
        n14418) );
  INVXL U35315 ( .A(weight_1[128]), .Y(n32710) );
  OAI22XL U35316 ( .A0(n32491), .A1(n32710), .B0(n32367), .B1(n16647), .Y(
        n14370) );
  INVXL U35317 ( .A(weight_1[146]), .Y(n32376) );
  OAI22XL U35318 ( .A0(n32491), .A1(n32368), .B0(n32376), .B1(n16647), .Y(
        n14372) );
  OAI22XL U35319 ( .A0(n32491), .A1(n32370), .B0(n32369), .B1(n16647), .Y(
        n14364) );
  OAI22XL U35320 ( .A0(n32491), .A1(n32371), .B0(n32378), .B1(n16647), .Y(
        n14349) );
  INVXL U35321 ( .A(weight_1[350]), .Y(n32404) );
  INVXL U35322 ( .A(weight_1[356]), .Y(n32717) );
  OAI22XL U35323 ( .A0(n32491), .A1(n32404), .B0(n32717), .B1(n16646), .Y(
        n14407) );
  INVXL U35324 ( .A(weight_1[374]), .Y(n32373) );
  INVXL U35325 ( .A(weight_1[380]), .Y(n32391) );
  OAI22XL U35326 ( .A0(n16645), .A1(n32373), .B0(n32391), .B1(n16646), .Y(
        n14411) );
  INVXL U35327 ( .A(weight_1[434]), .Y(n32389) );
  OAI22XL U35328 ( .A0(n16645), .A1(n32389), .B0(n32375), .B1(n16646), .Y(
        n14421) );
  OAI22XL U35329 ( .A0(n16650), .A1(n32379), .B0(n32372), .B1(n16646), .Y(
        n14424) );
  OAI22XL U35330 ( .A0(n32491), .A1(n32374), .B0(n32373), .B1(n16646), .Y(
        n14410) );
  OAI22XL U35331 ( .A0(n16650), .A1(n32375), .B0(n32380), .B1(n16646), .Y(
        n14422) );
  INVXL U35332 ( .A(weight_1[326]), .Y(n32392) );
  INVXL U35333 ( .A(weight_1[332]), .Y(n32400) );
  OAI22XL U35334 ( .A0(n16645), .A1(n32392), .B0(n32400), .B1(n16646), .Y(
        n14403) );
  INVXL U35335 ( .A(weight_1[152]), .Y(n32720) );
  OAI22XL U35336 ( .A0(n31071), .A1(n32376), .B0(n32720), .B1(n16647), .Y(
        n14373) );
  OAI22XL U35337 ( .A0(n32491), .A1(n32378), .B0(n32377), .B1(n16647), .Y(
        n14350) );
  OAI22XL U35338 ( .A0(n16650), .A1(n32380), .B0(n32379), .B1(n16646), .Y(
        n14423) );
  INVXL U35339 ( .A(weight_1[392]), .Y(n32397) );
  INVXL U35340 ( .A(weight_1[398]), .Y(n32734) );
  OAI22XL U35341 ( .A0(n16650), .A1(n32397), .B0(n32734), .B1(n16646), .Y(
        n14414) );
  INVXL U35342 ( .A(weight_1[400]), .Y(n32381) );
  OAI22XL U35343 ( .A0(n32491), .A1(n32452), .B0(n32381), .B1(n16646), .Y(
        n14252) );
  OAI22XL U35344 ( .A0(n31071), .A1(n32381), .B0(n32382), .B1(n16646), .Y(
        n14253) );
  INVXL U35345 ( .A(weight_1[412]), .Y(n32383) );
  OAI22XL U35346 ( .A0(n32491), .A1(n32382), .B0(n32383), .B1(n16646), .Y(
        n14254) );
  INVXL U35347 ( .A(weight_1[418]), .Y(n32752) );
  OAI22XL U35348 ( .A0(n31084), .A1(n32383), .B0(n32752), .B1(n16646), .Y(
        n14255) );
  INVXL U35349 ( .A(weight_1[436]), .Y(n32754) );
  OAI22XL U35350 ( .A0(n31071), .A1(n32754), .B0(n32384), .B1(n16646), .Y(
        n14259) );
  INVXL U35351 ( .A(weight_1[338]), .Y(n32399) );
  INVXL U35352 ( .A(weight_1[344]), .Y(n32405) );
  OAI22XL U35353 ( .A0(n16645), .A1(n32399), .B0(n32405), .B1(n16646), .Y(
        n14405) );
  OAI22XL U35354 ( .A0(n32491), .A1(n32385), .B0(n32386), .B1(n16646), .Y(
        n14261) );
  INVXL U35355 ( .A(weight_1[460]), .Y(n32756) );
  OAI22XL U35356 ( .A0(n16650), .A1(n32386), .B0(n32756), .B1(n16646), .Y(
        n14262) );
  OAI22XL U35357 ( .A0(n31077), .A1(n32759), .B0(n32387), .B1(n16646), .Y(
        n14266) );
  INVXL U35358 ( .A(weight_1[410]), .Y(n32396) );
  OAI22XL U35359 ( .A0(n32491), .A1(n32733), .B0(n32396), .B1(n16646), .Y(
        n14416) );
  OAI22XL U35360 ( .A0(n16645), .A1(n32388), .B0(n32401), .B1(n16646), .Y(
        n14268) );
  OAI22XL U35361 ( .A0(n16650), .A1(n32390), .B0(n32389), .B1(n16646), .Y(
        n14420) );
  OAI22XL U35362 ( .A0(n16645), .A1(n32391), .B0(n32398), .B1(n16646), .Y(
        n14412) );
  INVXL U35363 ( .A(weight_1[320]), .Y(n32721) );
  OAI22XL U35364 ( .A0(n32491), .A1(n32721), .B0(n32392), .B1(n16646), .Y(
        n14402) );
  OAI22XL U35365 ( .A0(n32491), .A1(n32394), .B0(n32393), .B1(n16647), .Y(
        n14366) );
  OAI22XL U35366 ( .A0(n32491), .A1(n32396), .B0(n32395), .B1(n16646), .Y(
        n14417) );
  OAI22XL U35367 ( .A0(n16645), .A1(n32398), .B0(n32397), .B1(n16646), .Y(
        n14413) );
  OAI22XL U35368 ( .A0(n16650), .A1(n32400), .B0(n32399), .B1(n16646), .Y(
        n14404) );
  OAI22XL U35369 ( .A0(n32491), .A1(n32463), .B0(n36145), .B1(n16646), .Y(
        n14348) );
  INVXL U35370 ( .A(weight_1[15]), .Y(n32403) );
  OAI22XL U35371 ( .A0(n32491), .A1(n32401), .B0(n32403), .B1(n16646), .Y(
        n14269) );
  INVXL U35372 ( .A(weight_1[363]), .Y(n32770) );
  INVXL U35373 ( .A(weight_1[369]), .Y(n32472) );
  OAI22XL U35374 ( .A0(n16645), .A1(n32770), .B0(n32472), .B1(n32777), .Y(
        n14328) );
  OAI22XL U35375 ( .A0(n16645), .A1(n32403), .B0(n32402), .B1(n16646), .Y(
        n14270) );
  OAI22XL U35376 ( .A0(n16650), .A1(n32405), .B0(n32404), .B1(n16646), .Y(
        n14406) );
  INVXL U35377 ( .A(weight_1[105]), .Y(n32761) );
  INVXL U35378 ( .A(weight_1[111]), .Y(n32406) );
  OAI22XL U35379 ( .A0(n32491), .A1(n32761), .B0(n32406), .B1(n32840), .Y(
        n14285) );
  INVXL U35380 ( .A(weight_1[117]), .Y(n32407) );
  OAI22XL U35381 ( .A0(n32491), .A1(n32406), .B0(n32407), .B1(n32840), .Y(
        n14286) );
  INVXL U35382 ( .A(weight_1[285]), .Y(n32715) );
  INVXL U35383 ( .A(weight_1[291]), .Y(n32762) );
  OAI22XL U35384 ( .A0(n31084), .A1(n32715), .B0(n32762), .B1(n32777), .Y(
        n14315) );
  INVXL U35385 ( .A(weight_1[36]), .Y(n32408) );
  INVXL U35386 ( .A(weight_1[42]), .Y(n32738) );
  OAI22XL U35387 ( .A0(n16650), .A1(n32408), .B0(n32738), .B1(n32840), .Y(
        n14517) );
  INVXL U35388 ( .A(weight_1[123]), .Y(n32413) );
  OAI22XL U35389 ( .A0(n32491), .A1(n32407), .B0(n32413), .B1(n32840), .Y(
        n14287) );
  INVXL U35390 ( .A(weight_1[30]), .Y(n32409) );
  OAI22XL U35391 ( .A0(n32491), .A1(n32409), .B0(n32408), .B1(n16648), .Y(
        n14516) );
  INVXL U35392 ( .A(weight_1[24]), .Y(n32410) );
  OAI22XL U35393 ( .A0(n16650), .A1(n32410), .B0(n32409), .B1(n26910), .Y(
        n14515) );
  OAI22XL U35394 ( .A0(n16650), .A1(n32411), .B0(n32410), .B1(n26910), .Y(
        n14514) );
  OAI22XL U35395 ( .A0(n31077), .A1(n32413), .B0(n32412), .B1(n32840), .Y(
        n14288) );
  OAI22XL U35396 ( .A0(n32491), .A1(n32414), .B0(n32724), .B1(n16648), .Y(
        n14511) );
  OAI22XL U35397 ( .A0(n16650), .A1(n32415), .B0(n36139), .B1(n16648), .Y(
        n14510) );
  INVXL U35398 ( .A(weight_1[475]), .Y(n32416) );
  OAI22XL U35399 ( .A0(n16645), .A1(n32416), .B0(n32415), .B1(n16648), .Y(
        n14509) );
  INVXL U35400 ( .A(weight_1[469]), .Y(n32417) );
  OAI22XL U35401 ( .A0(n16645), .A1(n32417), .B0(n32416), .B1(n16648), .Y(
        n14508) );
  INVXL U35402 ( .A(weight_1[463]), .Y(n32418) );
  OAI22XL U35403 ( .A0(n16645), .A1(n32418), .B0(n32417), .B1(n16648), .Y(
        n14507) );
  OAI22XL U35404 ( .A0(n31077), .A1(n32419), .B0(n32418), .B1(n16648), .Y(
        n14506) );
  INVXL U35405 ( .A(weight_1[87]), .Y(n32424) );
  INVXL U35406 ( .A(weight_1[93]), .Y(n32776) );
  OAI22XL U35407 ( .A0(n16650), .A1(n32424), .B0(n32776), .B1(n32840), .Y(
        n14282) );
  INVXL U35408 ( .A(weight_1[433]), .Y(n32420) );
  INVXL U35409 ( .A(weight_1[439]), .Y(n32728) );
  OAI22XL U35410 ( .A0(n16650), .A1(n32420), .B0(n32728), .B1(n16648), .Y(
        n14502) );
  OAI22XL U35411 ( .A0(n16650), .A1(n32421), .B0(n32420), .B1(n16648), .Y(
        n14501) );
  OAI22XL U35412 ( .A0(n16650), .A1(n32422), .B0(n32421), .B1(n16648), .Y(
        n14500) );
  OAI22XL U35413 ( .A0(n16650), .A1(n32423), .B0(n32422), .B1(n16648), .Y(
        n14499) );
  OAI22XL U35414 ( .A0(n32491), .A1(n32425), .B0(n32424), .B1(n32840), .Y(
        n14281) );
  INVXL U35415 ( .A(weight_1[141]), .Y(n32446) );
  OAI22XL U35416 ( .A0(n31084), .A1(n32446), .B0(n32426), .B1(n32840), .Y(
        n14291) );
  INVXL U35417 ( .A(weight_1[397]), .Y(n32698) );
  OAI22XL U35418 ( .A0(n16650), .A1(n32427), .B0(n32698), .B1(n16648), .Y(
        n14495) );
  OAI22XL U35419 ( .A0(n32491), .A1(n32428), .B0(n32427), .B1(n16648), .Y(
        n14494) );
  INVXL U35420 ( .A(weight_1[379]), .Y(n32429) );
  OAI22XL U35421 ( .A0(n32491), .A1(n32429), .B0(n32428), .B1(n16648), .Y(
        n14493) );
  INVXL U35422 ( .A(weight_1[373]), .Y(n32430) );
  OAI22XL U35423 ( .A0(n16645), .A1(n32430), .B0(n32429), .B1(n16648), .Y(
        n14492) );
  INVXL U35424 ( .A(weight_1[165]), .Y(n32718) );
  INVXL U35425 ( .A(weight_1[171]), .Y(n32692) );
  OAI22XL U35426 ( .A0(n32491), .A1(n32718), .B0(n32692), .B1(n32840), .Y(
        n14295) );
  INVXL U35427 ( .A(weight_1[367]), .Y(n32431) );
  OAI22XL U35428 ( .A0(n32491), .A1(n32431), .B0(n32430), .B1(n16648), .Y(
        n14491) );
  INVXL U35429 ( .A(weight_1[361]), .Y(n32434) );
  OAI22XL U35430 ( .A0(n16650), .A1(n32434), .B0(n32431), .B1(n16648), .Y(
        n14490) );
  INVXL U35431 ( .A(weight_1[63]), .Y(n32433) );
  OAI22XL U35432 ( .A0(n31084), .A1(n32433), .B0(n32432), .B1(n32840), .Y(
        n14278) );
  INVXL U35433 ( .A(weight_1[57]), .Y(n32437) );
  OAI22XL U35434 ( .A0(n32491), .A1(n32437), .B0(n32433), .B1(n16646), .Y(
        n14277) );
  INVXL U35435 ( .A(weight_1[355]), .Y(n32435) );
  OAI22XL U35436 ( .A0(n16650), .A1(n32435), .B0(n32434), .B1(n16648), .Y(
        n14489) );
  INVXL U35437 ( .A(weight_1[349]), .Y(n32436) );
  OAI22XL U35438 ( .A0(n16645), .A1(n32436), .B0(n32435), .B1(n16648), .Y(
        n14488) );
  INVXL U35439 ( .A(weight_1[343]), .Y(n32438) );
  OAI22XL U35440 ( .A0(n16650), .A1(n32438), .B0(n32436), .B1(n16648), .Y(
        n14487) );
  INVXL U35441 ( .A(weight_1[51]), .Y(n32442) );
  OAI22XL U35442 ( .A0(n32491), .A1(n32442), .B0(n32437), .B1(n16646), .Y(
        n14276) );
  INVXL U35443 ( .A(weight_1[337]), .Y(n32492) );
  OAI22XL U35444 ( .A0(n32491), .A1(n32492), .B0(n32438), .B1(n16648), .Y(
        n14486) );
  INVXL U35445 ( .A(weight_1[201]), .Y(n32439) );
  OAI22XL U35446 ( .A0(n16645), .A1(n32729), .B0(n32439), .B1(n32840), .Y(
        n14300) );
  INVXL U35447 ( .A(weight_1[207]), .Y(n32441) );
  OAI22XL U35448 ( .A0(n32491), .A1(n32439), .B0(n32441), .B1(n32840), .Y(
        n14301) );
  OAI22XL U35449 ( .A0(n16645), .A1(n32441), .B0(n32440), .B1(n32840), .Y(
        n14302) );
  INVXL U35450 ( .A(weight_1[45]), .Y(n32445) );
  OAI22XL U35451 ( .A0(n16650), .A1(n32445), .B0(n32442), .B1(n16646), .Y(
        n14275) );
  INVXL U35452 ( .A(weight_1[225]), .Y(n32699) );
  INVXL U35453 ( .A(weight_1[231]), .Y(n32691) );
  OAI22XL U35454 ( .A0(n16645), .A1(n32699), .B0(n32691), .B1(n32777), .Y(
        n14305) );
  INVXL U35455 ( .A(weight_1[243]), .Y(n32693) );
  INVXL U35456 ( .A(weight_1[249]), .Y(n32443) );
  OAI22XL U35457 ( .A0(n32491), .A1(n32693), .B0(n32443), .B1(n32777), .Y(
        n14308) );
  INVXL U35458 ( .A(weight_1[255]), .Y(n32444) );
  OAI22XL U35459 ( .A0(n16650), .A1(n32443), .B0(n32444), .B1(n32777), .Y(
        n14309) );
  INVXL U35460 ( .A(weight_1[261]), .Y(n32448) );
  OAI22XL U35461 ( .A0(n32491), .A1(n32444), .B0(n32448), .B1(n32777), .Y(
        n14310) );
  INVXL U35462 ( .A(weight_1[39]), .Y(n32773) );
  OAI22XL U35463 ( .A0(n16645), .A1(n32773), .B0(n32445), .B1(n16646), .Y(
        n14274) );
  OAI22XL U35464 ( .A0(n32491), .A1(n32447), .B0(n32446), .B1(n32840), .Y(
        n14290) );
  INVXL U35465 ( .A(weight_1[267]), .Y(n32705) );
  OAI22XL U35466 ( .A0(n16645), .A1(n32448), .B0(n32705), .B1(n32777), .Y(
        n14311) );
  INVXL U35467 ( .A(weight_1[235]), .Y(n32468) );
  INVXL U35468 ( .A(weight_1[241]), .Y(n32466) );
  OAI22XL U35469 ( .A0(n16645), .A1(n32468), .B0(n32466), .B1(n16646), .Y(
        n14469) );
  INVXL U35470 ( .A(weight_1[364]), .Y(n32453) );
  INVXL U35471 ( .A(weight_1[370]), .Y(n32449) );
  OAI22XL U35472 ( .A0(n31084), .A1(n32453), .B0(n32449), .B1(n16647), .Y(
        n14247) );
  INVXL U35473 ( .A(weight_1[346]), .Y(n32859) );
  INVXL U35474 ( .A(weight_1[352]), .Y(n32450) );
  OAI22XL U35475 ( .A0(n16645), .A1(n32859), .B0(n32450), .B1(n16647), .Y(
        n14244) );
  INVXL U35476 ( .A(weight_1[376]), .Y(n32451) );
  OAI22XL U35477 ( .A0(n32491), .A1(n32449), .B0(n32451), .B1(n16647), .Y(
        n14248) );
  INVXL U35478 ( .A(weight_1[358]), .Y(n32454) );
  OAI22XL U35479 ( .A0(n16645), .A1(n32450), .B0(n32454), .B1(n16647), .Y(
        n14245) );
  OAI22XL U35480 ( .A0(n16645), .A1(n32451), .B0(n32456), .B1(n16647), .Y(
        n14249) );
  INVXL U35481 ( .A(weight_1[388]), .Y(n32455) );
  OAI22XL U35482 ( .A0(n32491), .A1(n32455), .B0(n32452), .B1(n16647), .Y(
        n14251) );
  OAI22XL U35483 ( .A0(n31071), .A1(n32454), .B0(n32453), .B1(n16647), .Y(
        n14246) );
  OAI22XL U35484 ( .A0(n31077), .A1(n32456), .B0(n32455), .B1(n16647), .Y(
        n14250) );
  INVXL U35485 ( .A(conv_1[388]), .Y(n33146) );
  NAND4XL U35486 ( .A(conv_1[386]), .B(conv_1[387]), .C(n33089), .D(n33088), 
        .Y(n33148) );
  NAND3XL U35487 ( .A(n35463), .B(n33086), .C(n33093), .Y(n33147) );
  NAND2XL U35488 ( .A(n33148), .B(n33147), .Y(n32458) );
  NAND2XL U35489 ( .A(conv_1[388]), .B(n32458), .Y(n32457) );
  OAI211XL U35490 ( .A0(conv_1[388]), .A1(n32458), .B0(n33778), .C0(n32457), 
        .Y(n32459) );
  OAI211XL U35491 ( .A0(n35466), .A1(n33146), .B0(n34281), .C0(n32459), .Y(
        n16075) );
  INVXL U35492 ( .A(weight_1[145]), .Y(n32467) );
  INVXL U35493 ( .A(weight_1[151]), .Y(n32460) );
  INVXL U35494 ( .A(weight_1[223]), .Y(n32488) );
  INVXL U35495 ( .A(weight_1[229]), .Y(n32469) );
  INVXL U35496 ( .A(weight_1[157]), .Y(n32462) );
  INVXL U35497 ( .A(weight_1[175]), .Y(n32486) );
  INVXL U35498 ( .A(weight_1[181]), .Y(n32480) );
  INVXL U35499 ( .A(weight_1[187]), .Y(n32479) );
  INVXL U35500 ( .A(weight_1[247]), .Y(n32465) );
  INVXL U35501 ( .A(weight_1[253]), .Y(n32475) );
  INVXL U35502 ( .A(weight_1[163]), .Y(n32471) );
  INVXL U35503 ( .A(weight_1[259]), .Y(n32474) );
  INVXL U35504 ( .A(weight_1[265]), .Y(n32505) );
  INVXL U35505 ( .A(weight_1[139]), .Y(n32477) );
  INVXL U35506 ( .A(weight_1[199]), .Y(n32495) );
  INVXL U35507 ( .A(weight_1[205]), .Y(n32470) );
  INVXL U35508 ( .A(weight_1[211]), .Y(n32485) );
  INVXL U35509 ( .A(weight_1[169]), .Y(n32487) );
  INVXL U35510 ( .A(weight_1[375]), .Y(n32476) );
  INVXL U35511 ( .A(weight_1[381]), .Y(n32503) );
  INVXL U35512 ( .A(weight_1[133]), .Y(n32481) );
  INVXL U35513 ( .A(weight_1[441]), .Y(n32490) );
  INVXL U35514 ( .A(weight_1[217]), .Y(n32489) );
  INVXL U35515 ( .A(weight_1[331]), .Y(n32493) );
  INVXL U35516 ( .A(weight_1[325]), .Y(n32494) );
  INVXL U35517 ( .A(weight_1[319]), .Y(n32497) );
  INVXL U35518 ( .A(weight_1[313]), .Y(n32498) );
  INVXL U35519 ( .A(weight_1[283]), .Y(n32504) );
  INVXL U35520 ( .A(weight_1[289]), .Y(n32513) );
  INVXL U35521 ( .A(weight_1[307]), .Y(n32500) );
  INVXL U35522 ( .A(weight_1[411]), .Y(n32506) );
  INVXL U35523 ( .A(weight_1[417]), .Y(n32514) );
  INVXL U35524 ( .A(weight_1[429]), .Y(n32515) );
  INVXL U35525 ( .A(weight_1[301]), .Y(n32511) );
  INVXL U35526 ( .A(weight_1[387]), .Y(n32502) );
  INVXL U35527 ( .A(weight_1[277]), .Y(n32507) );
  INVXL U35528 ( .A(weight_1[271]), .Y(n32508) );
  INVXL U35529 ( .A(weight_1[295]), .Y(n32512) );
  INVXL U35530 ( .A(weight_1[423]), .Y(n32516) );
  OAI2BB1XL U35531 ( .A0N(conv_1[56]), .A1N(n32517), .B0(n35309), .Y(n32519)
         );
  INVXL U35532 ( .A(n32519), .Y(n32520) );
  OAI21XL U35533 ( .A0(n32521), .A1(n32520), .B0(n33822), .Y(n32523) );
  INVXL U35534 ( .A(conv_1[57]), .Y(n32522) );
  AOI32XL U35535 ( .A0(n35319), .A1(n32524), .A2(n32523), .B0(n32522), .B1(
        n32524), .Y(n16406) );
  AOI22XL U35536 ( .A0(n33712), .A1(n32526), .B0(conv_3[383]), .B1(n32623), 
        .Y(n32527) );
  NAND2XL U35537 ( .A(n32527), .B(n16649), .Y(n15490) );
  AOI22XL U35538 ( .A0(n32181), .A1(n32529), .B0(conv_3[324]), .B1(n33837), 
        .Y(n32530) );
  NAND2XL U35539 ( .A(n32530), .B(n16649), .Y(n15529) );
  ADDFX1 U35540 ( .A(conv_3[398]), .B(n33699), .CI(n32531), .CO(n32048), .S(
        n32533) );
  AOI22XL U35541 ( .A0(n30090), .A1(n32533), .B0(conv_3[398]), .B1(n32532), 
        .Y(n32534) );
  NAND2XL U35542 ( .A(n32534), .B(n16649), .Y(n15480) );
  NAND2BXL U35543 ( .AN(n32536), .B(n32535), .Y(n32538) );
  AOI211XL U35544 ( .A0(n32540), .A1(n32538), .B0(n36009), .C0(n32537), .Y(
        n32539) );
  NAND2XL U35545 ( .A(n32541), .B(n16649), .Y(n15539) );
  AOI22XL U35546 ( .A0(n33712), .A1(n32543), .B0(conv_3[66]), .B1(n32606), .Y(
        n32544) );
  NAND2XL U35547 ( .A(n32544), .B(n16649), .Y(n15702) );
  ADDFXL U35548 ( .A(conv_3[413]), .B(n32557), .CI(n32545), .CO(n32559), .S(
        n32547) );
  AOI22XL U35549 ( .A0(n33982), .A1(n32547), .B0(conv_3[413]), .B1(n32546), 
        .Y(n32548) );
  NAND2XL U35550 ( .A(n32548), .B(n16649), .Y(n15470) );
  AOI22XL U35551 ( .A0(n32660), .A1(n32550), .B0(conv_3[306]), .B1(n32614), 
        .Y(n32551) );
  NAND2XL U35552 ( .A(n32551), .B(n16649), .Y(n15542) );
  ADDFX1 U35553 ( .A(conv_3[71]), .B(n35599), .CI(n32552), .CO(n32164), .S(
        n32553) );
  AOI22XL U35554 ( .A0(n33712), .A1(n32553), .B0(conv_3[71]), .B1(n32606), .Y(
        n32554) );
  NAND2XL U35555 ( .A(n32554), .B(n16649), .Y(n15697) );
  INVXL U35556 ( .A(conv_3[415]), .Y(n32563) );
  AOI33XL U35557 ( .A0(conv_3[414]), .A1(n32559), .A2(n32558), .B0(n32557), 
        .B1(n32556), .B2(n32555), .Y(n32561) );
  AOI211XL U35558 ( .A0(n32563), .A1(n32561), .B0(n36042), .C0(n32560), .Y(
        n32562) );
  AOI2BB1XL U35559 ( .A0N(n32563), .A1N(n34227), .B0(n32562), .Y(n32564) );
  NAND2XL U35560 ( .A(n32564), .B(n16649), .Y(n15468) );
  AOI22XL U35561 ( .A0(n33778), .A1(n32567), .B0(conv_3[295]), .B1(n32566), 
        .Y(n32568) );
  NAND2XL U35562 ( .A(n32568), .B(n16649), .Y(n15548) );
  NAND2XL U35563 ( .A(n32574), .B(n16649), .Y(n15695) );
  OAI21XL U35564 ( .A0(n32578), .A1(n16655), .B0(n35778), .Y(n32577) );
  NAND2XL U35565 ( .A(n32580), .B(n16649), .Y(n15463) );
  AOI32XL U35566 ( .A0(conv_3[431]), .A1(n35775), .A2(n32582), .B0(n33790), 
        .B1(n32581), .Y(n32584) );
  AOI211XL U35567 ( .A0(n32586), .A1(n32584), .B0(n36042), .C0(n32583), .Y(
        n32585) );
  AOI2BB1XL U35568 ( .A0N(n32586), .A1N(n35778), .B0(n32585), .Y(n32587) );
  NAND2XL U35569 ( .A(n32587), .B(n16649), .Y(n15456) );
  INVXL U35570 ( .A(n32588), .Y(n32591) );
  AOI222XL U35571 ( .A0(conv_3[433]), .A1(n32591), .B0(conv_3[433]), .B1(
        n32590), .C0(n32589), .C1(n32588), .Y(n32592) );
  AOI22XL U35572 ( .A0(n32611), .A1(n32592), .B0(conv_3[433]), .B1(n33784), 
        .Y(n32593) );
  NAND2XL U35573 ( .A(n32593), .B(n16649), .Y(n15455) );
  AOI22XL U35574 ( .A0(n32656), .A1(n32595), .B0(conv_3[459]), .B1(n33774), 
        .Y(n32596) );
  NAND2XL U35575 ( .A(n32596), .B(n16649), .Y(n15439) );
  AOI32XL U35576 ( .A0(conv_3[281]), .A1(n32599), .A2(n32598), .B0(n32618), 
        .B1(n32597), .Y(n32601) );
  AOI211XL U35577 ( .A0(n32603), .A1(n32601), .B0(n36042), .C0(n32600), .Y(
        n32602) );
  AOI2BB1XL U35578 ( .A0N(n32603), .A1N(n34709), .B0(n32602), .Y(n32604) );
  NAND2XL U35579 ( .A(n32604), .B(n16649), .Y(n15556) );
  AOI22XL U35580 ( .A0(n33712), .A1(n32607), .B0(conv_3[65]), .B1(n32606), .Y(
        n32608) );
  NAND2XL U35581 ( .A(n32608), .B(n16649), .Y(n15703) );
  ADDFX1 U35582 ( .A(conv_3[311]), .B(n35732), .CI(n32609), .CO(n33111), .S(
        n32610) );
  AOI22XL U35583 ( .A0(n32611), .A1(n32610), .B0(conv_3[311]), .B1(n32614), 
        .Y(n32612) );
  NAND2XL U35584 ( .A(n32612), .B(n16649), .Y(n15537) );
  AOI22XL U35585 ( .A0(n32660), .A1(n32615), .B0(conv_3[310]), .B1(n32614), 
        .Y(n32616) );
  NAND2XL U35586 ( .A(n32616), .B(n16649), .Y(n15538) );
  AOI22XL U35587 ( .A0(n32656), .A1(n32620), .B0(conv_3[279]), .B1(n32619), 
        .Y(n32621) );
  NAND2XL U35588 ( .A(n32621), .B(n16649), .Y(n15559) );
  AOI22XL U35589 ( .A0(n33712), .A1(n32624), .B0(conv_3[381]), .B1(n32623), 
        .Y(n32625) );
  NAND2XL U35590 ( .A(n32625), .B(n16649), .Y(n15492) );
  OAI21XL U35591 ( .A0(n32629), .A1(n16654), .B0(n34227), .Y(n32628) );
  NAND2XL U35592 ( .A(n32631), .B(n16649), .Y(n15473) );
  ADDFX1 U35593 ( .A(conv_3[192]), .B(n32649), .CI(n32632), .CO(n32208), .S(
        n32633) );
  AOI22XL U35594 ( .A0(n32656), .A1(n32633), .B0(conv_3[192]), .B1(n32650), 
        .Y(n32634) );
  NAND2XL U35595 ( .A(n32634), .B(n16649), .Y(n15616) );
  INVXL U35596 ( .A(conv_3[115]), .Y(n32640) );
  NAND2XL U35597 ( .A(n34196), .B(n32636), .Y(n32635) );
  OAI21XL U35598 ( .A0(n34196), .A1(n32636), .B0(n32635), .Y(n32638) );
  AOI211XL U35599 ( .A0(n32640), .A1(n32638), .B0(n36009), .C0(n32637), .Y(
        n32639) );
  AOI2BB1XL U35600 ( .A0N(n32640), .A1N(n34200), .B0(n32639), .Y(n32641) );
  NAND2XL U35601 ( .A(n32641), .B(n16649), .Y(n15668) );
  INVXL U35602 ( .A(n32642), .Y(n32645) );
  AOI222XL U35603 ( .A0(conv_3[178]), .A1(n32645), .B0(conv_3[178]), .B1(
        n32644), .C0(n32643), .C1(n32642), .Y(n32646) );
  AOI22XL U35604 ( .A0(n16656), .A1(n32646), .B0(conv_3[178]), .B1(n35641), 
        .Y(n32647) );
  NAND2XL U35605 ( .A(n32647), .B(n16649), .Y(n15625) );
  AOI22XL U35606 ( .A0(n27932), .A1(n32651), .B0(conv_3[186]), .B1(n32650), 
        .Y(n32652) );
  NAND2XL U35607 ( .A(n32652), .B(n16649), .Y(n15622) );
  ADDFX1 U35608 ( .A(conv_3[114]), .B(n34196), .CI(n32653), .CO(n32636), .S(
        n32655) );
  AOI22XL U35609 ( .A0(n32656), .A1(n32655), .B0(conv_3[114]), .B1(n32654), 
        .Y(n32657) );
  NAND2XL U35610 ( .A(n32657), .B(n16649), .Y(n15669) );
  AOI22XL U35611 ( .A0(n32660), .A1(n32659), .B0(conv_3[173]), .B1(n35641), 
        .Y(n32661) );
  NAND2XL U35612 ( .A(n32661), .B(n16649), .Y(n15630) );
  AOI22XL U35613 ( .A0(n33712), .A1(n32663), .B0(conv_3[126]), .B1(n35572), 
        .Y(n32664) );
  NAND2XL U35614 ( .A(n32664), .B(n16649), .Y(n15662) );
  NAND2XL U35615 ( .A(n32670), .B(n16649), .Y(n15675) );
  NAND2XL U35616 ( .A(conv_2[89]), .B(n32675), .Y(n32674) );
  OAI22XL U35617 ( .A0(n32491), .A1(n32679), .B0(n32678), .B1(n26910), .Y(
        n14428) );
  OAI22XL U35618 ( .A0(n16645), .A1(n32681), .B0(n32680), .B1(n26910), .Y(
        n14437) );
  INVXL U35619 ( .A(weight_1[61]), .Y(n32684) );
  OAI22XL U35620 ( .A0(n32491), .A1(n32682), .B0(n32684), .B1(n26910), .Y(
        n14439) );
  OAI22XL U35621 ( .A0(n26906), .A1(n32684), .B0(n32683), .B1(n16647), .Y(
        n14440) );
  OAI22XL U35622 ( .A0(n32491), .A1(n32686), .B0(n32685), .B1(n16647), .Y(
        n14442) );
  ADDFX1 U35623 ( .A(conv_1[416]), .B(n35493), .CI(n32687), .CO(n34671), .S(
        n26522) );
  AOI22XL U35624 ( .A0(n33712), .A1(n32688), .B0(conv_1[417]), .B1(n35495), 
        .Y(n32689) );
  NAND2XL U35625 ( .A(n32689), .B(n34689), .Y(n16046) );
  INVXL U35626 ( .A(weight_1[206]), .Y(n32706) );
  INVXL U35627 ( .A(weight_1[212]), .Y(n32690) );
  OAI22XL U35628 ( .A0(n16650), .A1(n32706), .B0(n32690), .B1(n26910), .Y(
        n14383) );
  INVXL U35629 ( .A(weight_1[218]), .Y(n32747) );
  OAI22XL U35630 ( .A0(n32491), .A1(n32690), .B0(n32747), .B1(n26910), .Y(
        n14384) );
  INVXL U35631 ( .A(weight_1[237]), .Y(n32694) );
  OAI22XL U35632 ( .A0(n16645), .A1(n32691), .B0(n32694), .B1(n32777), .Y(
        n14306) );
  INVXL U35633 ( .A(weight_1[290]), .Y(n32725) );
  INVXL U35634 ( .A(weight_1[296]), .Y(n32707) );
  OAI22XL U35635 ( .A0(n32491), .A1(n32725), .B0(n32707), .B1(n16648), .Y(
        n14397) );
  INVXL U35636 ( .A(weight_1[278]), .Y(n32750) );
  INVXL U35637 ( .A(weight_1[284]), .Y(n32726) );
  OAI22XL U35638 ( .A0(n31071), .A1(n32750), .B0(n32726), .B1(n16646), .Y(
        n14395) );
  INVXL U35639 ( .A(weight_1[177]), .Y(n32695) );
  OAI22XL U35640 ( .A0(n31084), .A1(n32692), .B0(n32695), .B1(n32840), .Y(
        n14296) );
  OAI22XL U35641 ( .A0(n32491), .A1(n32694), .B0(n32693), .B1(n32777), .Y(
        n14307) );
  INVXL U35642 ( .A(weight_1[183]), .Y(n32702) );
  OAI22XL U35643 ( .A0(n16650), .A1(n32695), .B0(n32702), .B1(n32840), .Y(
        n14297) );
  INVXL U35644 ( .A(weight_1[403]), .Y(n32697) );
  OAI22XL U35645 ( .A0(n32491), .A1(n32697), .B0(n32696), .B1(n16648), .Y(
        n14497) );
  OAI22XL U35646 ( .A0(n16650), .A1(n32698), .B0(n32697), .B1(n16648), .Y(
        n14496) );
  OAI22XL U35647 ( .A0(n32491), .A1(n32700), .B0(n32699), .B1(n32777), .Y(
        n14304) );
  INVXL U35648 ( .A(weight_1[266]), .Y(n32701) );
  INVXL U35649 ( .A(weight_1[272]), .Y(n32751) );
  OAI22XL U35650 ( .A0(n32491), .A1(n32701), .B0(n32751), .B1(n16646), .Y(
        n14393) );
  INVXL U35651 ( .A(weight_1[260]), .Y(n32703) );
  OAI22XL U35652 ( .A0(n32491), .A1(n32703), .B0(n32701), .B1(n16646), .Y(
        n14392) );
  INVXL U35653 ( .A(weight_1[189]), .Y(n32730) );
  OAI22XL U35654 ( .A0(n16645), .A1(n32702), .B0(n32730), .B1(n32840), .Y(
        n14298) );
  INVXL U35655 ( .A(weight_1[254]), .Y(n32704) );
  OAI22XL U35656 ( .A0(n32491), .A1(n32704), .B0(n32703), .B1(n16648), .Y(
        n14391) );
  INVXL U35657 ( .A(weight_1[248]), .Y(n32714) );
  OAI22XL U35658 ( .A0(n16645), .A1(n32714), .B0(n32704), .B1(n32840), .Y(
        n14390) );
  INVXL U35659 ( .A(weight_1[273]), .Y(n32732) );
  OAI22XL U35660 ( .A0(n32491), .A1(n32705), .B0(n32732), .B1(n32777), .Y(
        n14312) );
  INVXL U35661 ( .A(weight_1[200]), .Y(n32742) );
  OAI22XL U35662 ( .A0(n32491), .A1(n32742), .B0(n32706), .B1(n32777), .Y(
        n14382) );
  INVXL U35663 ( .A(weight_1[302]), .Y(n32713) );
  OAI22XL U35664 ( .A0(n32491), .A1(n32707), .B0(n32713), .B1(n16647), .Y(
        n14398) );
  INVXL U35665 ( .A(weight_1[122]), .Y(n32711) );
  OAI22XL U35666 ( .A0(n16645), .A1(n32708), .B0(n32711), .B1(n16647), .Y(
        n14368) );
  INVXL U35667 ( .A(weight_1[159]), .Y(n32719) );
  OAI22XL U35668 ( .A0(n32491), .A1(n32709), .B0(n32719), .B1(n32840), .Y(
        n14293) );
  OAI22XL U35669 ( .A0(n31084), .A1(n32711), .B0(n32710), .B1(n16647), .Y(
        n14369) );
  OAI22XL U35670 ( .A0(n31084), .A1(n32713), .B0(n32712), .B1(n16648), .Y(
        n14399) );
  INVXL U35671 ( .A(weight_1[242]), .Y(n32741) );
  OAI22XL U35672 ( .A0(n32491), .A1(n32741), .B0(n32714), .B1(n26910), .Y(
        n14389) );
  INVXL U35673 ( .A(weight_1[279]), .Y(n32731) );
  OAI22XL U35674 ( .A0(n31084), .A1(n32731), .B0(n32715), .B1(n32777), .Y(
        n14314) );
  OAI22XL U35675 ( .A0(n16650), .A1(n32717), .B0(n32716), .B1(n16646), .Y(
        n14408) );
  OAI22XL U35676 ( .A0(n16650), .A1(n32719), .B0(n32718), .B1(n32840), .Y(
        n14294) );
  INVXL U35677 ( .A(weight_1[158]), .Y(n32735) );
  OAI22XL U35678 ( .A0(n16650), .A1(n32720), .B0(n32735), .B1(n26910), .Y(
        n14374) );
  OAI22XL U35679 ( .A0(n32491), .A1(n32722), .B0(n32721), .B1(n16646), .Y(
        n14401) );
  OAI22XL U35680 ( .A0(n32491), .A1(n32724), .B0(n32723), .B1(n26910), .Y(
        n14512) );
  OAI22XL U35681 ( .A0(n32491), .A1(n32726), .B0(n32725), .B1(n16646), .Y(
        n14396) );
  OAI22XL U35682 ( .A0(n32491), .A1(n32728), .B0(n32727), .B1(n16648), .Y(
        n14503) );
  OAI22XL U35683 ( .A0(n16650), .A1(n32730), .B0(n32729), .B1(n32840), .Y(
        n14299) );
  INVXL U35684 ( .A(weight_1[188]), .Y(n32745) );
  OAI22XL U35685 ( .A0(n16645), .A1(n32745), .B0(n32743), .B1(n16647), .Y(
        n14380) );
  OAI22XL U35686 ( .A0(n32491), .A1(n32732), .B0(n32731), .B1(n32777), .Y(
        n14313) );
  OAI22XL U35687 ( .A0(n32491), .A1(n32734), .B0(n32733), .B1(n16646), .Y(
        n14415) );
  INVXL U35688 ( .A(weight_1[164]), .Y(n32736) );
  OAI22XL U35689 ( .A0(n31071), .A1(n32735), .B0(n32736), .B1(n16648), .Y(
        n14375) );
  INVXL U35690 ( .A(weight_1[170]), .Y(n32739) );
  OAI22XL U35691 ( .A0(n31071), .A1(n32736), .B0(n32739), .B1(n26910), .Y(
        n14376) );
  OAI22XL U35692 ( .A0(n16650), .A1(n32738), .B0(n32737), .B1(n26910), .Y(
        n14518) );
  INVXL U35693 ( .A(weight_1[176]), .Y(n32740) );
  OAI22XL U35694 ( .A0(n31084), .A1(n32739), .B0(n32740), .B1(n16646), .Y(
        n14377) );
  INVXL U35695 ( .A(weight_1[182]), .Y(n32746) );
  OAI22XL U35696 ( .A0(n32491), .A1(n32740), .B0(n32746), .B1(n16646), .Y(
        n14378) );
  INVXL U35697 ( .A(weight_1[236]), .Y(n32744) );
  OAI22XL U35698 ( .A0(n32491), .A1(n32744), .B0(n32741), .B1(n16647), .Y(
        n14388) );
  OAI22XL U35699 ( .A0(n16650), .A1(n32743), .B0(n32742), .B1(n26910), .Y(
        n14381) );
  INVXL U35700 ( .A(weight_1[230]), .Y(n32748) );
  OAI22XL U35701 ( .A0(n32491), .A1(n32748), .B0(n32744), .B1(n16646), .Y(
        n14387) );
  OAI22XL U35702 ( .A0(n31077), .A1(n32746), .B0(n32745), .B1(n16647), .Y(
        n14379) );
  INVXL U35703 ( .A(weight_1[224]), .Y(n32749) );
  OAI22XL U35704 ( .A0(n31084), .A1(n32747), .B0(n32749), .B1(n26910), .Y(
        n14385) );
  INVXL U35705 ( .A(weight_1[315]), .Y(n32758) );
  INVXL U35706 ( .A(weight_1[321]), .Y(n32768) );
  OAI22XL U35707 ( .A0(n16650), .A1(n32758), .B0(n32768), .B1(n32777), .Y(
        n14320) );
  INVXL U35708 ( .A(weight_1[327]), .Y(n32767) );
  INVXL U35709 ( .A(weight_1[333]), .Y(n32769) );
  OAI22XL U35710 ( .A0(n16645), .A1(n32767), .B0(n32769), .B1(n32777), .Y(
        n14322) );
  OAI22XL U35711 ( .A0(n16645), .A1(n32752), .B0(n32753), .B1(n16646), .Y(
        n14256) );
  INVXL U35712 ( .A(weight_1[430]), .Y(n32755) );
  OAI22XL U35713 ( .A0(n31084), .A1(n32753), .B0(n32755), .B1(n16646), .Y(
        n14257) );
  OAI22XL U35714 ( .A0(n31077), .A1(n32755), .B0(n32754), .B1(n16646), .Y(
        n14258) );
  OAI22XL U35715 ( .A0(n32491), .A1(n32756), .B0(n32757), .B1(n16646), .Y(
        n14263) );
  OAI22XL U35716 ( .A0(n32491), .A1(n32757), .B0(n32760), .B1(n16646), .Y(
        n14264) );
  INVXL U35717 ( .A(weight_1[345]), .Y(n32771) );
  INVXL U35718 ( .A(weight_1[351]), .Y(n32779) );
  OAI22XL U35719 ( .A0(n31071), .A1(n32771), .B0(n32779), .B1(n32777), .Y(
        n14325) );
  INVXL U35720 ( .A(weight_1[309]), .Y(n32763) );
  OAI22XL U35721 ( .A0(n31084), .A1(n32763), .B0(n32758), .B1(n32777), .Y(
        n14319) );
  OAI22XL U35722 ( .A0(n32491), .A1(n32760), .B0(n32759), .B1(n16646), .Y(
        n14265) );
  INVXL U35723 ( .A(weight_1[99]), .Y(n32775) );
  OAI22XL U35724 ( .A0(n32491), .A1(n32775), .B0(n32761), .B1(n32840), .Y(
        n14284) );
  INVXL U35725 ( .A(weight_1[297]), .Y(n32765) );
  OAI22XL U35726 ( .A0(n16650), .A1(n32762), .B0(n32765), .B1(n32777), .Y(
        n14316) );
  INVXL U35727 ( .A(weight_1[303]), .Y(n32764) );
  OAI22XL U35728 ( .A0(n32491), .A1(n32764), .B0(n32763), .B1(n32777), .Y(
        n14318) );
  OAI22XL U35729 ( .A0(n16645), .A1(n32765), .B0(n32764), .B1(n32777), .Y(
        n14317) );
  INVXL U35730 ( .A(weight_1[33]), .Y(n32774) );
  OAI22XL U35731 ( .A0(n16650), .A1(n32766), .B0(n32774), .B1(n16646), .Y(
        n14272) );
  OAI22XL U35732 ( .A0(n16650), .A1(n32768), .B0(n32767), .B1(n32777), .Y(
        n14321) );
  INVXL U35733 ( .A(weight_1[339]), .Y(n32772) );
  OAI22XL U35734 ( .A0(n16650), .A1(n32769), .B0(n32772), .B1(n32777), .Y(
        n14323) );
  INVXL U35735 ( .A(weight_1[357]), .Y(n32778) );
  OAI22XL U35736 ( .A0(n16645), .A1(n32778), .B0(n32770), .B1(n32777), .Y(
        n14327) );
  OAI22XL U35737 ( .A0(n26906), .A1(n32772), .B0(n32771), .B1(n32777), .Y(
        n14324) );
  OAI22XL U35738 ( .A0(n32491), .A1(n32774), .B0(n32773), .B1(n16646), .Y(
        n14273) );
  OAI22XL U35739 ( .A0(n16645), .A1(n32776), .B0(n32775), .B1(n32840), .Y(
        n14283) );
  OAI22XL U35740 ( .A0(n32491), .A1(n32779), .B0(n32778), .B1(n32777), .Y(
        n14326) );
  OAI2BB1XL U35741 ( .A0N(conv_1[146]), .A1N(n34266), .B0(n32780), .Y(n32782)
         );
  AOI31XL U35742 ( .A0(n36020), .A1(n32781), .A2(n32782), .B0(n35549), .Y(
        n32787) );
  INVXL U35743 ( .A(n32782), .Y(n32783) );
  OAI21XL U35744 ( .A0(n32784), .A1(n32783), .B0(n33822), .Y(n32786) );
  INVXL U35745 ( .A(conv_1[147]), .Y(n32785) );
  AOI32XL U35746 ( .A0(n34271), .A1(n32787), .A2(n32786), .B0(n32785), .B1(
        n32787), .Y(n16316) );
  AOI32XL U35747 ( .A0(conv_3[146]), .A1(n32789), .A2(n33966), .B0(n33466), 
        .B1(n32788), .Y(n32791) );
  NAND2XL U35748 ( .A(n32793), .B(n32791), .Y(n32790) );
  OAI211XL U35749 ( .A0(n32793), .A1(n32791), .B0(n27932), .C0(n32790), .Y(
        n32792) );
  OAI211XL U35750 ( .A0(n34737), .A1(n32793), .B0(n16649), .C0(n32792), .Y(
        n15646) );
  NOR2BXL U35751 ( .AN(n32795), .B(n32794), .Y(n32797) );
  NAND2XL U35752 ( .A(conv_1[151]), .B(n32797), .Y(n32796) );
  OAI211XL U35753 ( .A0(conv_1[151]), .A1(n32797), .B0(n32656), .C0(n32796), 
        .Y(n32798) );
  OAI211XL U35754 ( .A0(n34048), .A1(n32799), .B0(n32798), .C0(n33067), .Y(
        n16312) );
  INVXL U35755 ( .A(weight_1[299]), .Y(n32809) );
  OAI22XL U35756 ( .A0(n16645), .A1(n32800), .B0(n32809), .B1(n26910), .Y(
        n14154) );
  INVXL U35757 ( .A(weight_1[263]), .Y(n32811) );
  OAI22XL U35758 ( .A0(n31084), .A1(n32801), .B0(n32811), .B1(n26910), .Y(
        n14148) );
  INVXL U35759 ( .A(weight_1[281]), .Y(n32805) );
  OAI22XL U35760 ( .A0(n31071), .A1(n32805), .B0(n32802), .B1(n16647), .Y(
        n14152) );
  INVXL U35761 ( .A(weight_1[269]), .Y(n32810) );
  INVXL U35762 ( .A(weight_1[275]), .Y(n32806) );
  OAI22XL U35763 ( .A0(n31077), .A1(n32810), .B0(n32806), .B1(n16647), .Y(
        n14150) );
  INVXL U35764 ( .A(weight_1[239]), .Y(n32803) );
  INVXL U35765 ( .A(weight_1[245]), .Y(n32808) );
  OAI22XL U35766 ( .A0(n16645), .A1(n32803), .B0(n32808), .B1(n26910), .Y(
        n14145) );
  INVXL U35767 ( .A(weight_1[233]), .Y(n32804) );
  OAI22XL U35768 ( .A0(n32967), .A1(n32804), .B0(n32803), .B1(n26910), .Y(
        n14144) );
  INVXL U35769 ( .A(weight_1[311]), .Y(n32812) );
  INVXL U35770 ( .A(weight_1[317]), .Y(n32814) );
  OAI22XL U35771 ( .A0(n31077), .A1(n32812), .B0(n32814), .B1(n16647), .Y(
        n14157) );
  INVXL U35772 ( .A(weight_1[227]), .Y(n32815) );
  OAI22XL U35773 ( .A0(n16645), .A1(n32815), .B0(n32804), .B1(n16647), .Y(
        n14143) );
  OAI22XL U35774 ( .A0(n32491), .A1(n32806), .B0(n32805), .B1(n26910), .Y(
        n14151) );
  OAI22XL U35775 ( .A0(n32491), .A1(n32808), .B0(n32807), .B1(n16647), .Y(
        n14146) );
  INVXL U35776 ( .A(weight_1[305]), .Y(n32813) );
  OAI22XL U35777 ( .A0(n32967), .A1(n32809), .B0(n32813), .B1(n26910), .Y(
        n14155) );
  OAI22XL U35778 ( .A0(n32491), .A1(n32811), .B0(n32810), .B1(n16647), .Y(
        n14149) );
  OAI22XL U35779 ( .A0(n16645), .A1(n32813), .B0(n32812), .B1(n26910), .Y(
        n14156) );
  INVXL U35780 ( .A(weight_1[323]), .Y(n32909) );
  OAI22XL U35781 ( .A0(n16650), .A1(n32814), .B0(n32909), .B1(n26910), .Y(
        n14158) );
  OAI22XL U35782 ( .A0(n31071), .A1(n32816), .B0(n32815), .B1(n16647), .Y(
        n14142) );
  INVXL U35783 ( .A(conv_1[106]), .Y(n32820) );
  NAND2XL U35784 ( .A(conv_1[106]), .B(n32818), .Y(n32817) );
  OAI211XL U35785 ( .A0(conv_1[106]), .A1(n32818), .B0(n32611), .C0(n32817), 
        .Y(n32819) );
  OAI211XL U35786 ( .A0(n35330), .A1(n32820), .B0(n32819), .C0(n33067), .Y(
        n16357) );
  INVXL U35787 ( .A(weight_1[112]), .Y(n32822) );
  INVXL U35788 ( .A(weight_1[118]), .Y(n32836) );
  OAI22XL U35789 ( .A0(n31084), .A1(n32822), .B0(n32836), .B1(n16648), .Y(
        n14205) );
  INVXL U35790 ( .A(weight_1[166]), .Y(n32824) );
  INVXL U35791 ( .A(weight_1[172]), .Y(n32823) );
  OAI22XL U35792 ( .A0(n16650), .A1(n32824), .B0(n32823), .B1(n16648), .Y(
        n14214) );
  INVXL U35793 ( .A(weight_1[184]), .Y(n32838) );
  INVXL U35794 ( .A(weight_1[190]), .Y(n32956) );
  OAI22XL U35795 ( .A0(n16650), .A1(n32838), .B0(n32956), .B1(n16648), .Y(
        n14217) );
  INVXL U35796 ( .A(weight_1[88]), .Y(n32833) );
  INVXL U35797 ( .A(weight_1[94]), .Y(n32821) );
  OAI22XL U35798 ( .A0(n16645), .A1(n32833), .B0(n32821), .B1(n16648), .Y(
        n14201) );
  INVXL U35799 ( .A(weight_1[100]), .Y(n32832) );
  OAI22XL U35800 ( .A0(n32967), .A1(n32821), .B0(n32832), .B1(n16648), .Y(
        n14202) );
  INVXL U35801 ( .A(weight_1[106]), .Y(n32831) );
  OAI22XL U35802 ( .A0(n16650), .A1(n32831), .B0(n32822), .B1(n16648), .Y(
        n14204) );
  INVXL U35803 ( .A(weight_1[178]), .Y(n32839) );
  OAI22XL U35804 ( .A0(n16650), .A1(n32823), .B0(n32839), .B1(n16648), .Y(
        n14215) );
  INVXL U35805 ( .A(weight_1[130]), .Y(n32834) );
  INVXL U35806 ( .A(weight_1[136]), .Y(n32830) );
  OAI22XL U35807 ( .A0(n16650), .A1(n32834), .B0(n32830), .B1(n16648), .Y(
        n14208) );
  INVXL U35808 ( .A(weight_1[160]), .Y(n32825) );
  OAI22XL U35809 ( .A0(n16650), .A1(n32825), .B0(n32824), .B1(n16648), .Y(
        n14213) );
  INVXL U35810 ( .A(weight_1[154]), .Y(n32826) );
  OAI22XL U35811 ( .A0(n16650), .A1(n32826), .B0(n32825), .B1(n16648), .Y(
        n14212) );
  INVXL U35812 ( .A(weight_1[148]), .Y(n32828) );
  OAI22XL U35813 ( .A0(n16650), .A1(n32828), .B0(n32826), .B1(n16648), .Y(
        n14211) );
  INVXL U35814 ( .A(weight_1[46]), .Y(n32827) );
  INVXL U35815 ( .A(weight_1[52]), .Y(n32843) );
  OAI22XL U35816 ( .A0(n32967), .A1(n32827), .B0(n32843), .B1(n16648), .Y(
        n14194) );
  INVXL U35817 ( .A(weight_1[40]), .Y(n32846) );
  OAI22XL U35818 ( .A0(n32967), .A1(n32846), .B0(n32827), .B1(n16648), .Y(
        n14193) );
  INVXL U35819 ( .A(weight_1[142]), .Y(n32829) );
  OAI22XL U35820 ( .A0(n16650), .A1(n32829), .B0(n32828), .B1(n16648), .Y(
        n14210) );
  OAI22XL U35821 ( .A0(n16650), .A1(n32830), .B0(n32829), .B1(n16648), .Y(
        n14209) );
  OAI22XL U35822 ( .A0(n16645), .A1(n32832), .B0(n32831), .B1(n16648), .Y(
        n14203) );
  INVXL U35823 ( .A(weight_1[82]), .Y(n32837) );
  OAI22XL U35824 ( .A0(n31084), .A1(n32837), .B0(n32833), .B1(n16648), .Y(
        n14200) );
  INVXL U35825 ( .A(weight_1[124]), .Y(n32835) );
  OAI22XL U35826 ( .A0(n32967), .A1(n32835), .B0(n32834), .B1(n16648), .Y(
        n14207) );
  OAI22XL U35827 ( .A0(n16650), .A1(n32836), .B0(n32835), .B1(n16648), .Y(
        n14206) );
  INVXL U35828 ( .A(weight_1[76]), .Y(n32841) );
  OAI22XL U35829 ( .A0(n16645), .A1(n32841), .B0(n32837), .B1(n16648), .Y(
        n14199) );
  OAI22XL U35830 ( .A0(n16650), .A1(n32839), .B0(n32838), .B1(n16648), .Y(
        n14216) );
  INVXL U35831 ( .A(weight_1[244]), .Y(n32968) );
  INVXL U35832 ( .A(weight_1[250]), .Y(n32849) );
  OAI22XL U35833 ( .A0(n16645), .A1(n32968), .B0(n32849), .B1(n32840), .Y(
        n14227) );
  INVXL U35834 ( .A(weight_1[64]), .Y(n32844) );
  INVXL U35835 ( .A(weight_1[70]), .Y(n32842) );
  OAI22XL U35836 ( .A0(n16650), .A1(n32844), .B0(n32842), .B1(n16648), .Y(
        n14197) );
  OAI22XL U35837 ( .A0(n31084), .A1(n32842), .B0(n32841), .B1(n16648), .Y(
        n14198) );
  INVXL U35838 ( .A(weight_1[58]), .Y(n32845) );
  OAI22XL U35839 ( .A0(n32967), .A1(n32843), .B0(n32845), .B1(n16648), .Y(
        n14195) );
  OAI22XL U35840 ( .A0(n16645), .A1(n32845), .B0(n32844), .B1(n16648), .Y(
        n14196) );
  INVXL U35841 ( .A(weight_1[34]), .Y(n32897) );
  OAI22XL U35842 ( .A0(n32967), .A1(n32897), .B0(n32846), .B1(n16648), .Y(
        n14192) );
  INVXL U35843 ( .A(weight_1[262]), .Y(n32850) );
  INVXL U35844 ( .A(weight_1[268]), .Y(n32853) );
  OAI22XL U35845 ( .A0(n16645), .A1(n32850), .B0(n32853), .B1(n16647), .Y(
        n14230) );
  INVXL U35846 ( .A(weight_1[274]), .Y(n32852) );
  INVXL U35847 ( .A(weight_1[280]), .Y(n32847) );
  OAI22XL U35848 ( .A0(n16645), .A1(n32852), .B0(n32847), .B1(n16647), .Y(
        n14232) );
  INVXL U35849 ( .A(weight_1[286]), .Y(n32848) );
  OAI22XL U35850 ( .A0(n16645), .A1(n32847), .B0(n32848), .B1(n16647), .Y(
        n14233) );
  INVXL U35851 ( .A(weight_1[292]), .Y(n32854) );
  OAI22XL U35852 ( .A0(n32967), .A1(n32848), .B0(n32854), .B1(n16647), .Y(
        n14234) );
  INVXL U35853 ( .A(weight_1[256]), .Y(n32851) );
  OAI22XL U35854 ( .A0(n16645), .A1(n32849), .B0(n32851), .B1(n16647), .Y(
        n14228) );
  OAI22XL U35855 ( .A0(n16645), .A1(n32851), .B0(n32850), .B1(n16647), .Y(
        n14229) );
  OAI22XL U35856 ( .A0(n16645), .A1(n32853), .B0(n32852), .B1(n16647), .Y(
        n14231) );
  INVXL U35857 ( .A(weight_1[298]), .Y(n32855) );
  OAI22XL U35858 ( .A0(n31071), .A1(n32854), .B0(n32855), .B1(n16647), .Y(
        n14235) );
  INVXL U35859 ( .A(weight_1[304]), .Y(n32863) );
  OAI22XL U35860 ( .A0(n31084), .A1(n32855), .B0(n32863), .B1(n16647), .Y(
        n14236) );
  INVXL U35861 ( .A(weight_1[328]), .Y(n32856) );
  INVXL U35862 ( .A(weight_1[334]), .Y(n32861) );
  OAI22XL U35863 ( .A0(n32967), .A1(n32856), .B0(n32861), .B1(n16647), .Y(
        n14241) );
  INVXL U35864 ( .A(weight_1[322]), .Y(n32857) );
  OAI22XL U35865 ( .A0(n32967), .A1(n32857), .B0(n32856), .B1(n16647), .Y(
        n14240) );
  INVXL U35866 ( .A(weight_1[310]), .Y(n32862) );
  INVXL U35867 ( .A(weight_1[316]), .Y(n32858) );
  OAI22XL U35868 ( .A0(n16645), .A1(n32862), .B0(n32858), .B1(n16647), .Y(
        n14238) );
  OAI22XL U35869 ( .A0(n16645), .A1(n32858), .B0(n32857), .B1(n16647), .Y(
        n14239) );
  INVXL U35870 ( .A(weight_1[340]), .Y(n32860) );
  OAI22XL U35871 ( .A0(n32967), .A1(n32860), .B0(n32859), .B1(n16647), .Y(
        n14243) );
  OAI22XL U35872 ( .A0(n16645), .A1(n32861), .B0(n32860), .B1(n16647), .Y(
        n14242) );
  OAI22XL U35873 ( .A0(n32491), .A1(n32863), .B0(n32862), .B1(n16647), .Y(
        n14237) );
  NAND2XL U35874 ( .A(n34028), .B(n32866), .Y(n32868) );
  OAI211XL U35875 ( .A0(n33432), .A1(n32869), .B0(n32868), .C0(n32867), .Y(
        n15935) );
  ADDFXL U35876 ( .A(conv_2[423]), .B(n32871), .CI(n32870), .CO(n28131), .S(
        n32872) );
  NAND2XL U35877 ( .A(n16657), .B(n32872), .Y(n32873) );
  OAI211XL U35878 ( .A0(n36053), .A1(n32874), .B0(n32873), .C0(n34105), .Y(
        n15247) );
  ADDFXL U35879 ( .A(conv_2[232]), .B(n32876), .CI(n32875), .CO(n29184), .S(
        n32877) );
  NAND2XL U35880 ( .A(n32611), .B(n32877), .Y(n32878) );
  OAI211XL U35881 ( .A0(n34458), .A1(n32879), .B0(n33815), .C0(n32878), .Y(
        n15051) );
  INVXL U35882 ( .A(conv_1[109]), .Y(n32885) );
  NOR2BXL U35883 ( .AN(n32881), .B(n32880), .Y(n32883) );
  NAND2XL U35884 ( .A(conv_1[109]), .B(n32883), .Y(n32882) );
  OAI211XL U35885 ( .A0(conv_1[109]), .A1(n32883), .B0(n33822), .C0(n32882), 
        .Y(n32884) );
  OAI211XL U35886 ( .A0(n35330), .A1(n32885), .B0(n35489), .C0(n32884), .Y(
        n16354) );
  ADDFX1 U35887 ( .A(conv_1[475]), .B(n32887), .CI(n32886), .CO(n29824), .S(
        n32888) );
  NAND2XL U35888 ( .A(n32656), .B(n32888), .Y(n32889) );
  OAI211XL U35889 ( .A0(n33506), .A1(n32890), .B0(n16652), .C0(n32889), .Y(
        n15988) );
  NAND2XL U35890 ( .A(n32656), .B(n32892), .Y(n32893) );
  OAI211XL U35891 ( .A0(n36053), .A1(n32894), .B0(n34669), .C0(n32893), .Y(
        n14918) );
  INVXL U35892 ( .A(weight_1[401]), .Y(n32895) );
  INVXL U35893 ( .A(weight_1[407]), .Y(n32908) );
  INVXL U35894 ( .A(weight_1[431]), .Y(n32917) );
  INVXL U35895 ( .A(weight_1[395]), .Y(n32896) );
  INVXL U35896 ( .A(weight_1[389]), .Y(n32899) );
  INVXL U35897 ( .A(weight_1[22]), .Y(n32911) );
  INVXL U35898 ( .A(weight_1[28]), .Y(n32898) );
  INVXL U35899 ( .A(weight_1[413]), .Y(n32907) );
  INVXL U35900 ( .A(weight_1[419]), .Y(n32916) );
  INVXL U35901 ( .A(weight_1[377]), .Y(n32938) );
  INVXL U35902 ( .A(weight_1[383]), .Y(n32900) );
  INVXL U35903 ( .A(weight_1[359]), .Y(n32903) );
  INVXL U35904 ( .A(weight_1[365]), .Y(n32940) );
  INVXL U35905 ( .A(weight_1[353]), .Y(n32904) );
  INVXL U35906 ( .A(weight_1[347]), .Y(n32945) );
  INVXL U35907 ( .A(weight_1[335]), .Y(n32948) );
  INVXL U35908 ( .A(weight_1[341]), .Y(n32946) );
  INVXL U35909 ( .A(weight_1[329]), .Y(n32949) );
  INVXL U35910 ( .A(weight_1[16]), .Y(n32965) );
  INVXL U35911 ( .A(weight_1[209]), .Y(n32913) );
  INVXL U35912 ( .A(weight_1[203]), .Y(n32914) );
  INVXL U35913 ( .A(weight_1[197]), .Y(n32915) );
  INVXL U35914 ( .A(weight_1[191]), .Y(n32919) );
  INVXL U35915 ( .A(weight_1[425]), .Y(n32918) );
  INVXL U35916 ( .A(weight_1[185]), .Y(n32920) );
  INVXL U35917 ( .A(weight_1[179]), .Y(n32963) );
  INVXL U35918 ( .A(weight_1[167]), .Y(n32924) );
  INVXL U35919 ( .A(weight_1[173]), .Y(n32964) );
  INVXL U35920 ( .A(weight_1[161]), .Y(n32925) );
  INVXL U35921 ( .A(weight_1[155]), .Y(n32926) );
  INVXL U35922 ( .A(weight_1[149]), .Y(n32927) );
  INVXL U35923 ( .A(weight_1[143]), .Y(n32928) );
  INVXL U35924 ( .A(weight_1[137]), .Y(n32931) );
  INVXL U35925 ( .A(weight_1[131]), .Y(n32932) );
  INVXL U35926 ( .A(weight_1[125]), .Y(n32933) );
  INVXL U35927 ( .A(weight_1[119]), .Y(n32934) );
  INVXL U35928 ( .A(weight_1[113]), .Y(n32935) );
  INVXL U35929 ( .A(weight_1[107]), .Y(n32936) );
  INVXL U35930 ( .A(weight_1[101]), .Y(n32937) );
  INVXL U35931 ( .A(weight_1[95]), .Y(n32941) );
  INVXL U35932 ( .A(weight_1[371]), .Y(n32939) );
  INVXL U35933 ( .A(weight_1[89]), .Y(n32942) );
  INVXL U35934 ( .A(weight_1[83]), .Y(n32943) );
  INVXL U35935 ( .A(weight_1[77]), .Y(n32944) );
  INVXL U35936 ( .A(weight_1[71]), .Y(n32947) );
  INVXL U35937 ( .A(weight_1[65]), .Y(n32950) );
  INVXL U35938 ( .A(weight_1[59]), .Y(n32951) );
  INVXL U35939 ( .A(weight_1[53]), .Y(n32952) );
  INVXL U35940 ( .A(weight_1[47]), .Y(n32953) );
  INVXL U35941 ( .A(weight_1[41]), .Y(n32954) );
  INVXL U35942 ( .A(weight_1[35]), .Y(n32955) );
  INVXL U35943 ( .A(weight_1[29]), .Y(n32957) );
  INVXL U35944 ( .A(weight_1[23]), .Y(n32958) );
  INVXL U35945 ( .A(weight_1[17]), .Y(n32960) );
  INVXL U35946 ( .A(weight_1[202]), .Y(n32973) );
  INVXL U35947 ( .A(weight_1[11]), .Y(n32961) );
  INVXL U35948 ( .A(weight_1[5]), .Y(n32962) );
  INVXL U35949 ( .A(weight_1[208]), .Y(n32972) );
  INVXL U35950 ( .A(weight_1[214]), .Y(n32975) );
  INVXL U35951 ( .A(weight_1[238]), .Y(n32969) );
  INVXL U35952 ( .A(weight_1[220]), .Y(n32974) );
  INVXL U35953 ( .A(weight_1[226]), .Y(n32971) );
  INVXL U35954 ( .A(weight_1[232]), .Y(n32970) );
  INVXL U35955 ( .A(conv_2[297]), .Y(n32981) );
  ADDFX1 U35956 ( .A(conv_2[296]), .B(n35957), .CI(n32976), .CO(n33136), .S(
        n30980) );
  NAND2XL U35957 ( .A(n35957), .B(n33136), .Y(n32977) );
  OAI21XL U35958 ( .A0(n35957), .A1(n33136), .B0(n32977), .Y(n32979) );
  AOI211XL U35959 ( .A0(n32981), .A1(n32979), .B0(n16655), .C0(n32978), .Y(
        n32980) );
  AOI2BB1XL U35960 ( .A0N(n32981), .A1N(n35963), .B0(n32980), .Y(n32982) );
  NAND2XL U35961 ( .A(n32982), .B(n34735), .Y(n15006) );
  ADDFXL U35962 ( .A(conv_2[258]), .B(n32984), .CI(n32983), .CO(n29409), .S(
        n32985) );
  NAND2XL U35963 ( .A(n16657), .B(n32985), .Y(n32986) );
  OAI211XL U35964 ( .A0(n34601), .A1(n32987), .B0(n32986), .C0(n34105), .Y(
        n15258) );
  NAND4XL U35965 ( .A(conv_1[191]), .B(conv_1[192]), .C(n32988), .D(n34085), 
        .Y(n34119) );
  INVXL U35966 ( .A(conv_1[192]), .Y(n34090) );
  NAND2XL U35967 ( .A(n32990), .B(n32989), .Y(n32991) );
  NAND3XL U35968 ( .A(n35365), .B(n34090), .C(n34086), .Y(n34118) );
  AOI22XL U35969 ( .A0(conv_1[193]), .A1(n34119), .B0(n34118), .B1(n34122), 
        .Y(n32993) );
  NAND2XL U35970 ( .A(conv_1[194]), .B(n32993), .Y(n32992) );
  OAI211XL U35971 ( .A0(conv_1[194]), .A1(n32993), .B0(n33778), .C0(n32992), 
        .Y(n32994) );
  OAI211XL U35972 ( .A0(n33853), .A1(n32995), .B0(n16652), .C0(n32994), .Y(
        n16269) );
  INVXL U35973 ( .A(conv_3[13]), .Y(n33153) );
  NAND4XL U35974 ( .A(conv_3[11]), .B(conv_3[12]), .C(n34378), .D(n32996), .Y(
        n33155) );
  NAND2XL U35975 ( .A(n34379), .B(n32997), .Y(n33154) );
  NAND2XL U35976 ( .A(n33155), .B(n33154), .Y(n32999) );
  NAND2XL U35977 ( .A(conv_3[13]), .B(n32999), .Y(n32998) );
  OAI211XL U35978 ( .A0(conv_3[13]), .A1(n32999), .B0(n33157), .C0(n32998), 
        .Y(n33000) );
  OAI211XL U35979 ( .A0(n34383), .A1(n33153), .B0(n33468), .C0(n33000), .Y(
        n15735) );
  ADDFXL U35980 ( .A(conv_3[20]), .B(n33002), .CI(n33001), .CO(n31274), .S(
        n33003) );
  NAND2XL U35981 ( .A(n16656), .B(n33003), .Y(n33004) );
  OAI211XL U35982 ( .A0(n35576), .A1(n33005), .B0(n16649), .C0(n33004), .Y(
        n15733) );
  INVXL U35983 ( .A(conv_3[266]), .Y(n33010) );
  OAI2BB1XL U35984 ( .A0N(n33006), .A1N(conv_3[264]), .B0(n33478), .Y(n35714)
         );
  OAI21XL U35985 ( .A0(conv_3[264]), .A1(n33007), .B0(n33480), .Y(n35712) );
  NAND2XL U35986 ( .A(n32611), .B(n33008), .Y(n33009) );
  OAI211XL U35987 ( .A0(n35713), .A1(n33010), .B0(n33468), .C0(n33009), .Y(
        n15567) );
  ADDFX1 U35988 ( .A(conv_3[473]), .B(n35810), .CI(n33011), .CO(n33015), .S(
        n33012) );
  NAND2XL U35989 ( .A(n24378), .B(n33012), .Y(n33013) );
  OAI211XL U35990 ( .A0(n35813), .A1(n33014), .B0(n16649), .C0(n33013), .Y(
        n15430) );
  ADDFX1 U35991 ( .A(conv_3[474]), .B(n35810), .CI(n33015), .CO(n32185), .S(
        n33016) );
  NAND2XL U35992 ( .A(n33822), .B(n33016), .Y(n33017) );
  OAI211XL U35993 ( .A0(n35813), .A1(n33018), .B0(n16649), .C0(n33017), .Y(
        n15429) );
  OAI21XL U35994 ( .A0(n33020), .A1(n33019), .B0(n33822), .Y(n33022) );
  AOI21XL U35995 ( .A0(n34742), .A1(n34438), .B0(conv_3[75]), .Y(n33021) );
  AOI32XL U35996 ( .A0(n35610), .A1(n34755), .A2(n33022), .B0(n33021), .B1(
        n34755), .Y(n15918) );
  INVXL U35997 ( .A(conv_3[272]), .Y(n33027) );
  NAND2XL U35998 ( .A(n24378), .B(n33025), .Y(n33026) );
  OAI211XL U35999 ( .A0(n34709), .A1(n33027), .B0(n33026), .C0(n35566), .Y(
        n15833) );
  INVXL U36000 ( .A(n33030), .Y(n33029) );
  OAI21XL U36001 ( .A0(n33029), .A1(n33028), .B0(n33157), .Y(n33033) );
  AOI31XL U36002 ( .A0(n36020), .A1(n33031), .A2(n33030), .B0(conv_1[211]), 
        .Y(n33032) );
  AOI32XL U36003 ( .A0(n35395), .A1(n33067), .A2(n33033), .B0(n33032), .B1(
        n33067), .Y(n16252) );
  AOI22XL U36004 ( .A0(conv_2[208]), .A1(n33036), .B0(n33035), .B1(n33034), 
        .Y(n33038) );
  NAND2XL U36005 ( .A(conv_2[209]), .B(n33038), .Y(n33037) );
  OAI211XL U36006 ( .A0(conv_2[209]), .A1(n33038), .B0(n30090), .C0(n33037), 
        .Y(n33039) );
  OAI211XL U36007 ( .A0(n34676), .A1(n33040), .B0(n35859), .C0(n33039), .Y(
        n15064) );
  AOI22XL U36008 ( .A0(conv_1[133]), .A1(n33043), .B0(n33042), .B1(n33041), 
        .Y(n33045) );
  NAND2XL U36009 ( .A(conv_1[134]), .B(n33045), .Y(n33044) );
  OAI211XL U36010 ( .A0(conv_1[134]), .A1(n33045), .B0(n32052), .C0(n33044), 
        .Y(n33046) );
  OAI211XL U36011 ( .A0(n34676), .A1(n33047), .B0(n34689), .C0(n33046), .Y(
        n16329) );
  AOI22XL U36012 ( .A0(conv_1[58]), .A1(n33050), .B0(n33049), .B1(n33048), .Y(
        n33052) );
  NAND2XL U36013 ( .A(conv_1[59]), .B(n33052), .Y(n33051) );
  OAI211XL U36014 ( .A0(conv_1[59]), .A1(n33052), .B0(n32611), .C0(n33051), 
        .Y(n33053) );
  OAI211XL U36015 ( .A0(n34676), .A1(n33054), .B0(n16652), .C0(n33053), .Y(
        n16404) );
  OAI21XL U36016 ( .A0(n33056), .A1(n33055), .B0(n32660), .Y(n33060) );
  AOI31XL U36017 ( .A0(n36020), .A1(n33058), .A2(n33057), .B0(conv_2[302]), 
        .Y(n33059) );
  AOI32XL U36018 ( .A0(n35976), .A1(n34621), .A2(n33060), .B0(n33059), .B1(
        n34621), .Y(n15291) );
  INVXL U36019 ( .A(n33063), .Y(n33062) );
  OAI21XL U36020 ( .A0(n33062), .A1(n33061), .B0(n32181), .Y(n33066) );
  AOI31XL U36021 ( .A0(n36020), .A1(n33064), .A2(n33063), .B0(conv_1[166]), 
        .Y(n33065) );
  AOI32XL U36022 ( .A0(n35346), .A1(n33067), .A2(n33066), .B0(n33065), .B1(
        n33067), .Y(n16297) );
  NAND2XL U36023 ( .A(n33554), .B(n33068), .Y(n33074) );
  XOR2XL U36024 ( .A(DP_OP_5168J1_124_9881_n12), .B(affine_1[9]), .Y(n33071)
         );
  XOR2X1 U36025 ( .A(n33072), .B(n33071), .Y(n33073) );
  INVXL U36026 ( .A(n33075), .Y(n33561) );
  NAND4XL U36027 ( .A(conv_2[326]), .B(conv_2[327]), .C(n33079), .D(n33933), 
        .Y(n33233) );
  INVXL U36028 ( .A(conv_2[327]), .Y(n33938) );
  NAND2XL U36029 ( .A(n33081), .B(n33080), .Y(n33082) );
  NAND2XL U36030 ( .A(n35982), .B(n33082), .Y(n33934) );
  NAND3XL U36031 ( .A(n35982), .B(n33938), .C(n33934), .Y(n33232) );
  NAND2XL U36032 ( .A(n33233), .B(n33232), .Y(n33084) );
  NAND2XL U36033 ( .A(conv_2[328]), .B(n33084), .Y(n33083) );
  OAI211XL U36034 ( .A0(conv_2[328]), .A1(n33084), .B0(n32181), .C0(n33083), 
        .Y(n33085) );
  OAI211XL U36035 ( .A0(n35986), .A1(n33231), .B0(n34735), .C0(n33085), .Y(
        n14985) );
  AOI32XL U36036 ( .A0(n33089), .A1(n33088), .A2(n33087), .B0(n33086), .B1(
        n35463), .Y(n33091) );
  NAND2XL U36037 ( .A(n33093), .B(n33091), .Y(n33090) );
  OAI211XL U36038 ( .A0(n33093), .A1(n33091), .B0(n33778), .C0(n33090), .Y(
        n33092) );
  OAI211XL U36039 ( .A0(n35466), .A1(n33093), .B0(n34544), .C0(n33092), .Y(
        n16076) );
  OAI32XL U36040 ( .A0(conv_2[238]), .A1(n33097), .A2(n33096), .B0(n33095), 
        .B1(n33094), .Y(n33099) );
  NAND2XL U36041 ( .A(conv_2[239]), .B(n33099), .Y(n33098) );
  OAI211XL U36042 ( .A0(conv_2[239]), .A1(n33099), .B0(n32052), .C0(n33098), 
        .Y(n33100) );
  OAI211XL U36043 ( .A0(n33853), .A1(n33101), .B0(n35859), .C0(n33100), .Y(
        n15044) );
  AOI22XL U36044 ( .A0(conv_2[58]), .A1(n33104), .B0(n33103), .B1(n33102), .Y(
        n33106) );
  NAND2XL U36045 ( .A(conv_2[59]), .B(n33106), .Y(n33105) );
  OAI211XL U36046 ( .A0(conv_2[59]), .A1(n33106), .B0(n16657), .C0(n33105), 
        .Y(n33107) );
  OAI211XL U36047 ( .A0(n34520), .A1(n33108), .B0(n33815), .C0(n33107), .Y(
        n15164) );
  NAND3XL U36048 ( .A(conv_3[312]), .B(n33111), .C(n33109), .Y(n34031) );
  NAND3BXL U36049 ( .AN(n33111), .B(n35732), .C(n33110), .Y(n34030) );
  INVXL U36050 ( .A(conv_3[313]), .Y(n34034) );
  AOI22XL U36051 ( .A0(conv_3[313]), .A1(n34031), .B0(n34030), .B1(n34034), 
        .Y(n33113) );
  NAND2XL U36052 ( .A(conv_3[314]), .B(n33113), .Y(n33112) );
  OAI211XL U36053 ( .A0(conv_3[314]), .A1(n33113), .B0(n16656), .C0(n33112), 
        .Y(n33114) );
  OAI211XL U36054 ( .A0(n34789), .A1(n33115), .B0(n33468), .C0(n33114), .Y(
        n15534) );
  AOI22XL U36055 ( .A0(conv_1[208]), .A1(n33118), .B0(n33117), .B1(n33116), 
        .Y(n33120) );
  NAND2XL U36056 ( .A(conv_1[209]), .B(n33120), .Y(n33119) );
  OAI211XL U36057 ( .A0(conv_1[209]), .A1(n33120), .B0(n24378), .C0(n33119), 
        .Y(n33121) );
  OAI211XL U36058 ( .A0(n33853), .A1(n33122), .B0(n34689), .C0(n33121), .Y(
        n16254) );
  NAND2XL U36059 ( .A(n33251), .B(n35289), .Y(n33250) );
  INVXL U36060 ( .A(conv_1[43]), .Y(n33253) );
  OAI32XL U36061 ( .A0(conv_1[43]), .A1(n33251), .A2(n35289), .B0(n33250), 
        .B1(n33253), .Y(n33125) );
  NAND2XL U36062 ( .A(conv_1[44]), .B(n33125), .Y(n33124) );
  OAI211XL U36063 ( .A0(conv_1[44]), .A1(n33125), .B0(n16657), .C0(n33124), 
        .Y(n33126) );
  OAI211XL U36064 ( .A0(n34676), .A1(n33127), .B0(n34689), .C0(n33126), .Y(
        n16419) );
  OAI211XL U36065 ( .A0(conv_1[374]), .A1(n33132), .B0(n33982), .C0(n33131), 
        .Y(n33133) );
  INVXL U36066 ( .A(conv_2[298]), .Y(n33294) );
  NAND3XL U36067 ( .A(conv_2[297]), .B(n33136), .C(n33135), .Y(n33296) );
  OR3XL U36068 ( .A(n33136), .B(conv_2[297]), .C(n33135), .Y(n33295) );
  NAND2XL U36069 ( .A(n33296), .B(n33295), .Y(n33138) );
  NAND2XL U36070 ( .A(conv_2[298]), .B(n33138), .Y(n33137) );
  OAI211XL U36071 ( .A0(conv_2[298]), .A1(n33138), .B0(n28751), .C0(n33137), 
        .Y(n33139) );
  OAI211XL U36072 ( .A0(n35963), .A1(n33294), .B0(n34735), .C0(n33139), .Y(
        n15005) );
  INVXL U36073 ( .A(conv_2[403]), .Y(n33256) );
  NAND4XL U36074 ( .A(conv_2[401]), .B(conv_2[402]), .C(n33953), .D(n36033), 
        .Y(n33258) );
  OAI21XL U36075 ( .A0(conv_2[400]), .A1(n33142), .B0(n34634), .Y(n36032) );
  INVXL U36076 ( .A(conv_2[402]), .Y(n33957) );
  NAND3XL U36077 ( .A(n36034), .B(n34634), .C(n33957), .Y(n33257) );
  NAND2XL U36078 ( .A(n33258), .B(n33257), .Y(n33144) );
  NAND2XL U36079 ( .A(conv_2[403]), .B(n33144), .Y(n33143) );
  OAI211XL U36080 ( .A0(conv_2[403]), .A1(n33144), .B0(n16657), .C0(n33143), 
        .Y(n33145) );
  OAI211XL U36081 ( .A0(n36031), .A1(n33256), .B0(n35859), .C0(n33145), .Y(
        n14935) );
  OAI211XL U36082 ( .A0(conv_1[389]), .A1(n33150), .B0(n32181), .C0(n33149), 
        .Y(n33151) );
  NAND2XL U36083 ( .A(conv_3[14]), .B(n33158), .Y(n33156) );
  NAND2XL U36084 ( .A(n32611), .B(n33161), .Y(n33165) );
  OAI21XL U36085 ( .A0(n33166), .A1(n33162), .B0(n33157), .Y(n33163) );
  OAI2BB1XL U36086 ( .A0N(n33506), .A1N(n33163), .B0(conv_1[470]), .Y(n33164)
         );
  OAI211XL U36087 ( .A0(n33166), .A1(n33165), .B0(n16652), .C0(n33164), .Y(
        n15993) );
  OAI2BB1XL U36088 ( .A0N(conv_2[506]), .A1N(n33704), .B0(n36081), .Y(n33170)
         );
  AOI31XL U36089 ( .A0(n36020), .A1(n33705), .A2(n33170), .B0(n16651), .Y(
        n33175) );
  INVXL U36090 ( .A(n33170), .Y(n33171) );
  OAI21XL U36091 ( .A0(n33172), .A1(n33171), .B0(n32181), .Y(n33174) );
  AOI32XL U36092 ( .A0(n36091), .A1(n33175), .A2(n33174), .B0(n33173), .B1(
        n33175), .Y(n14866) );
  NAND2XL U36093 ( .A(n24378), .B(n33176), .Y(n33180) );
  OAI21XL U36094 ( .A0(n33181), .A1(n33177), .B0(n33982), .Y(n33178) );
  OAI2BB1XL U36095 ( .A0N(n35466), .A1N(n33178), .B0(conv_1[380]), .Y(n33179)
         );
  OAI211XL U36096 ( .A0(n33181), .A1(n33180), .B0(n16652), .C0(n33179), .Y(
        n16083) );
  NAND2XL U36097 ( .A(n32656), .B(n33182), .Y(n33186) );
  OAI21XL U36098 ( .A0(n33187), .A1(n33183), .B0(n33788), .Y(n33184) );
  OAI2BB1XL U36099 ( .A0N(n35408), .A1N(n33184), .B0(conv_1[230]), .Y(n33185)
         );
  OAI211XL U36100 ( .A0(n33187), .A1(n33186), .B0(n34682), .C0(n33185), .Y(
        n16233) );
  NAND2XL U36101 ( .A(n31735), .B(n33188), .Y(n33192) );
  OAI21XL U36102 ( .A0(n33189), .A1(n33193), .B0(n16657), .Y(n33190) );
  OAI2BB1XL U36103 ( .A0N(n35368), .A1N(n33190), .B0(conv_1[185]), .Y(n33191)
         );
  OAI211XL U36104 ( .A0(n33193), .A1(n33192), .B0(n16652), .C0(n33191), .Y(
        n16278) );
  NAND2XL U36105 ( .A(n24378), .B(n33194), .Y(n33198) );
  OAI21XL U36106 ( .A0(n33195), .A1(n33199), .B0(n16657), .Y(n33196) );
  OAI2BB1XL U36107 ( .A0N(n35945), .A1N(n33196), .B0(conv_2[250]), .Y(n33197)
         );
  OAI211XL U36108 ( .A0(n33199), .A1(n33198), .B0(n35859), .C0(n33197), .Y(
        n15038) );
  OR4XL U36109 ( .A(n33202), .B(n33201), .C(n33200), .D(n35275), .Y(n33438) );
  NAND2XL U36110 ( .A(n35275), .B(n33203), .Y(n33437) );
  NAND2XL U36111 ( .A(n33438), .B(n33437), .Y(n33205) );
  NAND2XL U36112 ( .A(conv_1[28]), .B(n33205), .Y(n33204) );
  OAI211XL U36113 ( .A0(conv_1[28]), .A1(n33205), .B0(n33778), .C0(n33204), 
        .Y(n33206) );
  OAI211XL U36114 ( .A0(n35278), .A1(n33436), .B0(n34544), .C0(n33206), .Y(
        n16435) );
  OR4XL U36115 ( .A(n33209), .B(n33208), .C(n33207), .D(n35541), .Y(n33354) );
  NAND2XL U36116 ( .A(n35541), .B(n33210), .Y(n33353) );
  NAND2XL U36117 ( .A(n33354), .B(n33353), .Y(n33212) );
  NAND2XL U36118 ( .A(conv_1[493]), .B(n33212), .Y(n33211) );
  OAI211XL U36119 ( .A0(conv_1[493]), .A1(n33212), .B0(n34666), .C0(n33211), 
        .Y(n33213) );
  OAI211XL U36120 ( .A0(n35544), .A1(n33352), .B0(n16652), .C0(n33213), .Y(
        n15970) );
  NAND2XL U36121 ( .A(n24378), .B(n33214), .Y(n33218) );
  OAI21XL U36122 ( .A0(n33219), .A1(n33215), .B0(n24499), .Y(n33216) );
  OAI2BB1XL U36123 ( .A0N(n34080), .A1N(n33216), .B0(conv_1[259]), .Y(n33217)
         );
  OAI211XL U36124 ( .A0(n33219), .A1(n33218), .B0(n33217), .C0(n35489), .Y(
        n16204) );
  OAI21XL U36125 ( .A0(n33699), .A1(n33696), .B0(n33697), .Y(n33224) );
  NAND2XL U36126 ( .A(n33698), .B(n33224), .Y(n33223) );
  OAI211XL U36127 ( .A0(n33698), .A1(n33224), .B0(n32181), .C0(n33223), .Y(
        n33225) );
  OAI211XL U36128 ( .A0(n33703), .A1(n33698), .B0(n16649), .C0(n33225), .Y(
        n15476) );
  ADDFX1 U36129 ( .A(conv_3[266]), .B(n33480), .CI(n33226), .CO(n33481), .S(
        n33008) );
  AOI21XL U36130 ( .A0(n33481), .A1(n33480), .B0(n33227), .Y(n33229) );
  NAND2XL U36131 ( .A(conv_3[267]), .B(n33229), .Y(n33228) );
  OAI211XL U36132 ( .A0(conv_3[267]), .A1(n33229), .B0(n24378), .C0(n33228), 
        .Y(n33230) );
  OAI211XL U36133 ( .A0(n35713), .A1(n33479), .B0(n16649), .C0(n33230), .Y(
        n15566) );
  AOI22XL U36134 ( .A0(conv_2[328]), .A1(n33233), .B0(n33232), .B1(n33231), 
        .Y(n33235) );
  NAND2XL U36135 ( .A(conv_2[329]), .B(n33235), .Y(n33234) );
  OAI211XL U36136 ( .A0(conv_2[329]), .A1(n33235), .B0(n30090), .C0(n33234), 
        .Y(n33236) );
  OAI211XL U36137 ( .A0(n33442), .A1(n33237), .B0(n35859), .C0(n33236), .Y(
        n14984) );
  OAI21XL U36138 ( .A0(n36001), .A1(n33241), .B0(n35330), .Y(n33240) );
  NAND2XL U36139 ( .A(n33243), .B(n34696), .Y(n16345) );
  NAND2XL U36140 ( .A(n33245), .B(n33244), .Y(n33247) );
  OAI21XL U36141 ( .A0(n36009), .A1(n33247), .B0(n33506), .Y(n33246) );
  AOI32XL U36142 ( .A0(n32660), .A1(n33248), .A2(n33247), .B0(conv_1[478]), 
        .B1(n33246), .Y(n33249) );
  NAND2XL U36143 ( .A(n33249), .B(n34281), .Y(n15985) );
  AOI22XL U36144 ( .A0(conv_2[403]), .A1(n33258), .B0(n33257), .B1(n33256), 
        .Y(n33260) );
  NAND2XL U36145 ( .A(conv_2[404]), .B(n33260), .Y(n33259) );
  OAI211XL U36146 ( .A0(conv_2[404]), .A1(n33260), .B0(n33788), .C0(n33259), 
        .Y(n33261) );
  OAI211XL U36147 ( .A0(n34676), .A1(n33262), .B0(n33815), .C0(n33261), .Y(
        n14934) );
  NAND2XL U36148 ( .A(n33264), .B(n33263), .Y(n33266) );
  OAI21XL U36149 ( .A0(n36009), .A1(n33266), .B0(n35934), .Y(n33265) );
  AOI32XL U36150 ( .A0(n34028), .A1(n33267), .A2(n33266), .B0(conv_2[223]), 
        .B1(n33265), .Y(n33268) );
  NAND2XL U36151 ( .A(n33268), .B(n34735), .Y(n15055) );
  NAND4XL U36152 ( .A(conv_1[401]), .B(conv_1[402]), .C(n35471), .D(n35479), 
        .Y(n34692) );
  NAND3XL U36153 ( .A(n35480), .B(n33654), .C(n33269), .Y(n34691) );
  AOI22XL U36154 ( .A0(conv_1[403]), .A1(n34692), .B0(n34691), .B1(n34695), 
        .Y(n33271) );
  NAND2XL U36155 ( .A(conv_1[404]), .B(n33271), .Y(n33270) );
  OAI211XL U36156 ( .A0(conv_1[404]), .A1(n33271), .B0(n32052), .C0(n33270), 
        .Y(n33272) );
  OAI211XL U36157 ( .A0(n33442), .A1(n33273), .B0(n34696), .C0(n33272), .Y(
        n16059) );
  NAND2XL U36158 ( .A(n33275), .B(n33274), .Y(n33277) );
  OAI21XL U36159 ( .A0(n34389), .A1(n33277), .B0(n34177), .Y(n33276) );
  AOI32XL U36160 ( .A0(n30090), .A1(n33278), .A2(n33277), .B0(conv_2[478]), 
        .B1(n33276), .Y(n33279) );
  NAND2XL U36161 ( .A(n33279), .B(n34735), .Y(n14885) );
  NAND4XL U36162 ( .A(conv_3[326]), .B(conv_3[327]), .C(n33281), .D(n33280), 
        .Y(n34067) );
  NAND3XL U36163 ( .A(n33283), .B(n33842), .C(n33282), .Y(n34066) );
  INVXL U36164 ( .A(conv_3[328]), .Y(n34070) );
  AOI22XL U36165 ( .A0(conv_3[328]), .A1(n34067), .B0(n34066), .B1(n34070), 
        .Y(n33285) );
  NAND2XL U36166 ( .A(conv_3[329]), .B(n33285), .Y(n33284) );
  OAI211XL U36167 ( .A0(conv_3[329]), .A1(n33285), .B0(n28751), .C0(n33284), 
        .Y(n33286) );
  OAI211XL U36168 ( .A0(n34789), .A1(n33287), .B0(n33468), .C0(n33286), .Y(
        n15524) );
  NAND2XL U36169 ( .A(n33289), .B(n33288), .Y(n33291) );
  OAI21XL U36170 ( .A0(n36042), .A1(n33291), .B0(n34447), .Y(n33290) );
  NAND2XL U36171 ( .A(n33293), .B(n34735), .Y(n15135) );
  NAND2XL U36172 ( .A(conv_2[299]), .B(n33298), .Y(n33297) );
  OAI211XL U36173 ( .A0(conv_2[299]), .A1(n33298), .B0(n30090), .C0(n33297), 
        .Y(n33299) );
  NAND2XL U36174 ( .A(n33302), .B(n33301), .Y(n33305) );
  OAI21XL U36175 ( .A0(n16655), .A1(n33305), .B0(n33303), .Y(n33304) );
  NAND2XL U36176 ( .A(n33307), .B(n35588), .Y(n15395) );
  NAND2XL U36177 ( .A(n33309), .B(n33308), .Y(n33311) );
  OAI21XL U36178 ( .A0(n36009), .A1(n33311), .B0(n35826), .Y(n33310) );
  AOI32XL U36179 ( .A0(n33822), .A1(n33312), .A2(n33311), .B0(conv_3[493]), 
        .B1(n33310), .Y(n33313) );
  NAND2XL U36180 ( .A(n33313), .B(n35588), .Y(n15415) );
  INVXL U36181 ( .A(conv_3[237]), .Y(n33880) );
  NAND2XL U36182 ( .A(n33315), .B(n33314), .Y(n33316) );
  AOI32XL U36183 ( .A0(conv_3[236]), .A1(n33879), .A2(n33877), .B0(n35673), 
        .B1(n33879), .Y(n33318) );
  NAND2XL U36184 ( .A(n33880), .B(n33318), .Y(n33317) );
  OAI211XL U36185 ( .A0(n33880), .A1(n33318), .B0(n33822), .C0(n33317), .Y(
        n33319) );
  OAI211XL U36186 ( .A0(n35676), .A1(n33880), .B0(n16649), .C0(n33319), .Y(
        n15586) );
  NAND3XL U36187 ( .A(conv_2[417]), .B(n36044), .C(n33321), .Y(n34037) );
  AOI21XL U36188 ( .A0(n36045), .A1(n36044), .B0(conv_2[417]), .Y(n36049) );
  NAND2XL U36189 ( .A(n36045), .B(n36049), .Y(n34036) );
  INVXL U36190 ( .A(conv_2[418]), .Y(n34040) );
  AOI22XL U36191 ( .A0(conv_2[418]), .A1(n34037), .B0(n34036), .B1(n34040), 
        .Y(n33323) );
  NAND2XL U36192 ( .A(conv_2[419]), .B(n33323), .Y(n33322) );
  OAI211XL U36193 ( .A0(conv_2[419]), .A1(n33323), .B0(n32656), .C0(n33322), 
        .Y(n33324) );
  OAI211XL U36194 ( .A0(n34789), .A1(n33325), .B0(n34735), .C0(n33324), .Y(
        n14924) );
  INVXL U36195 ( .A(n33328), .Y(n33327) );
  AOI221XL U36196 ( .A0(n33327), .A1(n16656), .B0(n33326), .B1(n16656), .C0(
        n33714), .Y(n33331) );
  AOI31XL U36197 ( .A0(n36020), .A1(n33329), .A2(n33328), .B0(conv_3[526]), 
        .Y(n33330) );
  OAI21XL U36198 ( .A0(n33331), .A1(n33330), .B0(n33550), .Y(n15852) );
  ADDFXL U36199 ( .A(affine_2[45]), .B(affine_2[46]), .CI(n33336), .CO(n33337), 
        .S(n33333) );
  ADDFX1 U36200 ( .A(n33344), .B(n33343), .CI(n33342), .CO(n33345), .S(n28401)
         );
  ADDFXL U36201 ( .A(affine_2[29]), .B(affine_2[30]), .CI(n33346), .CO(n33347), 
        .S(n33343) );
  AOI22XL U36202 ( .A0(conv_1[493]), .A1(n33354), .B0(n33353), .B1(n33352), 
        .Y(n33356) );
  NAND2XL U36203 ( .A(conv_1[494]), .B(n33356), .Y(n33355) );
  OAI211XL U36204 ( .A0(conv_1[494]), .A1(n33356), .B0(n34666), .C0(n33355), 
        .Y(n33357) );
  OAI211XL U36205 ( .A0(n33442), .A1(n33358), .B0(n16652), .C0(n33357), .Y(
        n15969) );
  ADDFXL U36206 ( .A(affine_2[13]), .B(affine_2[14]), .CI(n33363), .CO(n33364), 
        .S(n33360) );
  AOI221XL U36207 ( .A0(n33371), .A1(n24499), .B0(n33370), .B1(n16656), .C0(
        n33624), .Y(n33376) );
  OAI211XL U36208 ( .A0(n33629), .A1(n33373), .B0(n32052), .C0(n33372), .Y(
        n33374) );
  OAI211XL U36209 ( .A0(n33376), .A1(n33375), .B0(n33815), .C0(n33374), .Y(
        n14848) );
  INVXL U36210 ( .A(n33379), .Y(n33378) );
  AOI221XL U36211 ( .A0(n33378), .A1(n24378), .B0(n33377), .B1(n16657), .C0(
        n33687), .Y(n33383) );
  AOI31XL U36212 ( .A0(n36020), .A1(n33380), .A2(n33379), .B0(n16651), .Y(
        n33381) );
  OAI21XL U36213 ( .A0(n33383), .A1(n33382), .B0(n33381), .Y(n14933) );
  AOI221XL U36214 ( .A0(n33385), .A1(n34028), .B0(n33384), .B1(n16656), .C0(
        n35495), .Y(n33390) );
  INVXL U36215 ( .A(conv_1[414]), .Y(n33389) );
  OAI211XL U36216 ( .A0(n35493), .A1(n33387), .B0(n33822), .C0(n33386), .Y(
        n33388) );
  OAI211XL U36217 ( .A0(n33390), .A1(n33389), .B0(n34682), .C0(n33388), .Y(
        n16049) );
  AOI221XL U36218 ( .A0(n33392), .A1(n36020), .B0(n33391), .B1(n16656), .C0(
        n35510), .Y(n33397) );
  INVXL U36219 ( .A(conv_1[429]), .Y(n33396) );
  OAI211XL U36220 ( .A0(intadd_1_B_2_), .A1(n33394), .B0(n32181), .C0(n33393), 
        .Y(n33395) );
  OAI211XL U36221 ( .A0(n33397), .A1(n33396), .B0(n16652), .C0(n33395), .Y(
        n16034) );
  INVXL U36222 ( .A(n33539), .Y(n33541) );
  OAI21XL U36223 ( .A0(n33403), .A1(n35499), .B0(n33402), .Y(n33540) );
  NAND2XL U36224 ( .A(conv_1[422]), .B(n33540), .Y(n33538) );
  NAND2XL U36225 ( .A(n33541), .B(n33538), .Y(intadd_1_CI) );
  NAND2XL U36226 ( .A(n33554), .B(n33404), .Y(n33410) );
  XOR2X1 U36227 ( .A(n33406), .B(DP_OP_5166J1_122_9881_n13), .Y(n33408) );
  XOR2XL U36228 ( .A(DP_OP_5166J1_122_9881_n12), .B(affine_1[29]), .Y(n33407)
         );
  AOI221XL U36229 ( .A0(n33415), .A1(n36020), .B0(n33414), .B1(n16656), .C0(
        n34531), .Y(n33420) );
  INVXL U36230 ( .A(conv_2[381]), .Y(n33419) );
  OAI211XL U36231 ( .A0(n34529), .A1(n33417), .B0(n33788), .C0(n33416), .Y(
        n33418) );
  OAI211XL U36232 ( .A0(n33420), .A1(n33419), .B0(n34669), .C0(n33418), .Y(
        n14952) );
  OAI21XL U36233 ( .A0(n33422), .A1(n33421), .B0(n33157), .Y(n33426) );
  AOI21XL U36234 ( .A0(n34769), .A1(n33424), .B0(conv_1[495]), .Y(n33425) );
  AOI32XL U36235 ( .A0(n33427), .A1(n34773), .A2(n33426), .B0(n33425), .B1(
        n34773), .Y(n15968) );
  OAI21XL U36236 ( .A0(n33429), .A1(n33428), .B0(n33157), .Y(n33431) );
  AOI21XL U36237 ( .A0(n34769), .A1(n34498), .B0(conv_1[525]), .Y(n33430) );
  AOI32XL U36238 ( .A0(n33432), .A1(n34773), .A2(n33431), .B0(n33430), .B1(
        n34773), .Y(n15938) );
  OAI21XL U36239 ( .A0(n33988), .A1(n33433), .B0(n32181), .Y(n33435) );
  AOI21XL U36240 ( .A0(n34769), .A1(n33990), .B0(conv_1[30]), .Y(n33434) );
  AOI32XL U36241 ( .A0(n35302), .A1(n34773), .A2(n33435), .B0(n33434), .B1(
        n34773), .Y(n16433) );
  OAI211XL U36242 ( .A0(conv_1[29]), .A1(n33440), .B0(n33778), .C0(n33439), 
        .Y(n33441) );
  AOI221XL U36243 ( .A0(n33446), .A1(n16656), .B0(n33445), .B1(n16656), .C0(
        n33444), .Y(n33452) );
  INVXL U36244 ( .A(conv_3[37]), .Y(n33451) );
  OAI211XL U36245 ( .A0(n33449), .A1(n33448), .B0(n33778), .C0(n33447), .Y(
        n33450) );
  OAI211XL U36246 ( .A0(n33452), .A1(n33451), .B0(n16649), .C0(n33450), .Y(
        n15721) );
  AOI221XL U36247 ( .A0(n33455), .A1(n16656), .B0(n33454), .B1(n16656), .C0(
        n33453), .Y(n33460) );
  OAI211XL U36248 ( .A0(n35914), .A1(n33457), .B0(n28751), .C0(n33456), .Y(
        n33458) );
  OAI211XL U36249 ( .A0(n33460), .A1(n33459), .B0(n35859), .C0(n33458), .Y(
        n15078) );
  AOI221XL U36250 ( .A0(n33463), .A1(n16656), .B0(n33462), .B1(n16656), .C0(
        n33461), .Y(n33470) );
  OAI211XL U36251 ( .A0(n33466), .A1(n33465), .B0(n36020), .C0(n33464), .Y(
        n33467) );
  OAI211XL U36252 ( .A0(n33470), .A1(n33469), .B0(n33468), .C0(n33467), .Y(
        n15648) );
  AOI221XL U36253 ( .A0(n33472), .A1(n36020), .B0(n33471), .B1(n16656), .C0(
        n33747), .Y(n33477) );
  OAI211XL U36254 ( .A0(n33752), .A1(n33474), .B0(n16656), .C0(n33473), .Y(
        n33475) );
  OAI211XL U36255 ( .A0(n33477), .A1(n33476), .B0(n16649), .C0(n33475), .Y(
        n15508) );
  NAND3XL U36256 ( .A(conv_3[267]), .B(n33481), .C(n33478), .Y(n33907) );
  NAND3BXL U36257 ( .AN(n33481), .B(n33480), .C(n33479), .Y(n33906) );
  NAND2XL U36258 ( .A(n33907), .B(n33906), .Y(n33483) );
  NAND2XL U36259 ( .A(conv_3[268]), .B(n33483), .Y(n33482) );
  OAI211XL U36260 ( .A0(conv_3[268]), .A1(n33483), .B0(n16657), .C0(n33482), 
        .Y(n33484) );
  OAI211XL U36261 ( .A0(n35713), .A1(n33905), .B0(n33468), .C0(n33484), .Y(
        n15565) );
  NAND4XL U36262 ( .A(conv_1[236]), .B(conv_1[237]), .C(n34276), .D(n34275), 
        .Y(n33848) );
  INVXL U36263 ( .A(conv_1[237]), .Y(n34280) );
  NAND3XL U36264 ( .A(n34274), .B(n35404), .C(n34280), .Y(n33847) );
  NAND2XL U36265 ( .A(n33848), .B(n33847), .Y(n33486) );
  OAI21XL U36266 ( .A0(n36042), .A1(n33486), .B0(n35408), .Y(n33485) );
  NAND2XL U36267 ( .A(n33487), .B(n16652), .Y(n16225) );
  OAI21XL U36268 ( .A0(n33488), .A1(n36042), .B0(n35327), .Y(n33489) );
  AOI32XL U36269 ( .A0(n34769), .A1(n33489), .A2(n34699), .B0(conv_1[60]), 
        .B1(n33489), .Y(n33490) );
  NAND2XL U36270 ( .A(n34773), .B(n33490), .Y(n16403) );
  AOI32XL U36271 ( .A0(n34769), .A1(n33492), .A2(n34493), .B0(conv_1[120]), 
        .B1(n33492), .Y(n33493) );
  NAND2XL U36272 ( .A(n34773), .B(n33493), .Y(n16343) );
  OAI21XL U36273 ( .A0(n33494), .A1(n36042), .B0(n34057), .Y(n33495) );
  AOI32XL U36274 ( .A0(n34769), .A1(n33495), .A2(n34438), .B0(conv_1[75]), 
        .B1(n33495), .Y(n33496) );
  NAND2XL U36275 ( .A(n34773), .B(n33496), .Y(n16388) );
  INVXL U36276 ( .A(conv_1[165]), .Y(n33499) );
  OAI21XL U36277 ( .A0(n33497), .A1(n36042), .B0(n35346), .Y(n33498) );
  AOI32XL U36278 ( .A0(n34769), .A1(n33499), .A2(n34433), .B0(conv_1[165]), 
        .B1(n33498), .Y(n33500) );
  NAND2XL U36279 ( .A(n33500), .B(n34773), .Y(n16298) );
  INVXL U36280 ( .A(conv_1[135]), .Y(n33504) );
  OAI21XL U36281 ( .A0(n33502), .A1(n16655), .B0(n34271), .Y(n33503) );
  AOI32XL U36282 ( .A0(n34769), .A1(n33504), .A2(n34740), .B0(conv_1[135]), 
        .B1(n33503), .Y(n33505) );
  NAND2XL U36283 ( .A(n33505), .B(n34773), .Y(n16328) );
  OAI21XL U36284 ( .A0(n33507), .A1(n36042), .B0(n33506), .Y(n33508) );
  AOI32XL U36285 ( .A0(n34769), .A1(n33510), .A2(n33509), .B0(conv_1[465]), 
        .B1(n33508), .Y(n33511) );
  NAND2XL U36286 ( .A(n33511), .B(n34773), .Y(n15998) );
  OAI21XL U36287 ( .A0(n33512), .A1(n16655), .B0(n35319), .Y(n33513) );
  AOI32XL U36288 ( .A0(n34769), .A1(n33514), .A2(n34507), .B0(conv_1[45]), 
        .B1(n33513), .Y(n33515) );
  NAND2XL U36289 ( .A(n33515), .B(n34773), .Y(n16418) );
  INVXL U36290 ( .A(conv_1[285]), .Y(n33518) );
  AOI32XL U36291 ( .A0(n33516), .A1(n34325), .A2(n34455), .B0(n16655), .B1(
        n34325), .Y(n33517) );
  AOI32XL U36292 ( .A0(n34769), .A1(n33518), .A2(n34455), .B0(conv_1[285]), 
        .B1(n33517), .Y(n33519) );
  NAND2XL U36293 ( .A(n33519), .B(n34773), .Y(n16178) );
  AOI32XL U36294 ( .A0(n33520), .A1(n35487), .A2(n34229), .B0(n16655), .B1(
        n35487), .Y(n33521) );
  AOI32XL U36295 ( .A0(n34769), .A1(n33522), .A2(n34229), .B0(conv_1[405]), 
        .B1(n33521), .Y(n33523) );
  NAND2XL U36296 ( .A(n33523), .B(n34773), .Y(n16058) );
  OAI2BB1XL U36297 ( .A0N(n36020), .A1N(n33524), .B0(n34080), .Y(n33525) );
  AOI32XL U36298 ( .A0(n34769), .A1(n33526), .A2(n34422), .B0(conv_1[255]), 
        .B1(n33525), .Y(n33527) );
  NAND2XL U36299 ( .A(n33527), .B(n34773), .Y(n16208) );
  INVXL U36300 ( .A(conv_1[480]), .Y(n33531) );
  OAI2BB1XL U36301 ( .A0N(n36020), .A1N(n33528), .B0(n35544), .Y(n33529) );
  AOI32XL U36302 ( .A0(n34769), .A1(n33531), .A2(n33530), .B0(conv_1[480]), 
        .B1(n33529), .Y(n33532) );
  NAND2XL U36303 ( .A(n33532), .B(n34773), .Y(n15983) );
  AOI32XL U36304 ( .A0(n33533), .A1(n35417), .A2(n33535), .B0(n16654), .B1(
        n35417), .Y(n33534) );
  AOI32XL U36305 ( .A0(n34769), .A1(n33536), .A2(n33535), .B0(conv_1[240]), 
        .B1(n33534), .Y(n33537) );
  NAND2XL U36306 ( .A(n33537), .B(n34773), .Y(n16223) );
  AOI221XL U36307 ( .A0(n33539), .A1(n32656), .B0(n33538), .B1(n33982), .C0(
        n35510), .Y(n33544) );
  OAI21XL U36308 ( .A0(n33544), .A1(n33543), .B0(n33542), .Y(n16041) );
  AOI221XL U36309 ( .A0(n33547), .A1(n34028), .B0(n33546), .B1(n16657), .C0(
        n33545), .Y(n33552) );
  AOI31XL U36310 ( .A0(n16657), .A1(n33549), .A2(n33548), .B0(conv_3[241]), 
        .Y(n33551) );
  OAI21XL U36311 ( .A0(n33552), .A1(n33551), .B0(n33550), .Y(n15871) );
  NAND2XL U36312 ( .A(n33554), .B(n33553), .Y(n33560) );
  ADDFX1 U36313 ( .A(DP_OP_5167J1_123_9881_n16), .B(DP_OP_5167J1_123_9881_n14), 
        .CI(n33555), .CO(n33556), .S(n25244) );
  XOR2X1 U36314 ( .A(n33556), .B(DP_OP_5167J1_123_9881_n13), .Y(n33558) );
  XOR2XL U36315 ( .A(DP_OP_5167J1_123_9881_n12), .B(affine_1[19]), .Y(n33557)
         );
  NAND2XL U36316 ( .A(n33565), .B(n33564), .Y(n16482) );
  AOI221XL U36317 ( .A0(n33568), .A1(n36020), .B0(n33567), .B1(n16656), .C0(
        n33566), .Y(n33574) );
  INVXL U36318 ( .A(conv_2[8]), .Y(n33573) );
  OAI211XL U36319 ( .A0(n33571), .A1(n33570), .B0(n36020), .C0(n33569), .Y(
        n33572) );
  OAI211XL U36320 ( .A0(n33574), .A1(n33573), .B0(n35859), .C0(n33572), .Y(
        n15200) );
  AOI221XL U36321 ( .A0(n33577), .A1(n30090), .B0(n33576), .B1(n31735), .C0(
        n33575), .Y(n33583) );
  INVXL U36322 ( .A(conv_2[516]), .Y(n33582) );
  OAI211XL U36323 ( .A0(n33580), .A1(n33579), .B0(n16657), .C0(n33578), .Y(
        n33581) );
  OAI211XL U36324 ( .A0(n33583), .A1(n33582), .B0(n34669), .C0(n33581), .Y(
        n14862) );
  AOI221XL U36325 ( .A0(n33585), .A1(n33982), .B0(n33584), .B1(n33912), .C0(
        n33986), .Y(n33591) );
  OAI211XL U36326 ( .A0(n33588), .A1(n33587), .B0(n16657), .C0(n33586), .Y(
        n33589) );
  OAI211XL U36327 ( .A0(n33591), .A1(n33590), .B0(n34669), .C0(n33589), .Y(
        n15178) );
  AOI221XL U36328 ( .A0(n33592), .A1(n33788), .B0(n33594), .B1(n33712), .C0(
        n33986), .Y(n33597) );
  NAND3BXL U36329 ( .AN(n33594), .B(n33593), .C(n33982), .Y(n33595) );
  OAI211XL U36330 ( .A0(n33597), .A1(n33596), .B0(n33815), .C0(n33595), .Y(
        n15183) );
  AOI221XL U36331 ( .A0(n33600), .A1(n33778), .B0(n33599), .B1(n16657), .C0(
        n33598), .Y(n33605) );
  INVXL U36332 ( .A(conv_2[486]), .Y(n33604) );
  OAI211XL U36333 ( .A0(n34132), .A1(n33602), .B0(n16656), .C0(n33601), .Y(
        n33603) );
  OAI211XL U36334 ( .A0(n33605), .A1(n33604), .B0(n34669), .C0(n33603), .Y(
        n14882) );
  AOI221XL U36335 ( .A0(n33608), .A1(n33157), .B0(n33607), .B1(n24499), .C0(
        n33606), .Y(n33614) );
  INVXL U36336 ( .A(conv_2[460]), .Y(n33613) );
  OAI211XL U36337 ( .A0(n33611), .A1(n33610), .B0(n16656), .C0(n33609), .Y(
        n33612) );
  OAI211XL U36338 ( .A0(n33614), .A1(n33613), .B0(n34669), .C0(n33612), .Y(
        n14898) );
  AOI221XL U36339 ( .A0(n33617), .A1(n32660), .B0(n33616), .B1(n33912), .C0(
        n33615), .Y(n33623) );
  OAI211XL U36340 ( .A0(n33620), .A1(n33619), .B0(n33822), .C0(n33618), .Y(
        n33621) );
  OAI211XL U36341 ( .A0(n33623), .A1(n33622), .B0(n35859), .C0(n33621), .Y(
        n15190) );
  AOI221XL U36342 ( .A0(n33626), .A1(n33982), .B0(n33625), .B1(n33912), .C0(
        n33624), .Y(n33632) );
  INVXL U36343 ( .A(conv_2[533]), .Y(n33631) );
  OAI211XL U36344 ( .A0(n33629), .A1(n33628), .B0(n30090), .C0(n33627), .Y(
        n33630) );
  OAI211XL U36345 ( .A0(n33632), .A1(n33631), .B0(n35859), .C0(n33630), .Y(
        n14850) );
  AOI221XL U36346 ( .A0(n33635), .A1(n33778), .B0(n33634), .B1(n16657), .C0(
        n33633), .Y(n33641) );
  OAI211XL U36347 ( .A0(n33638), .A1(n33637), .B0(n33157), .C0(n33636), .Y(
        n33639) );
  OAI211XL U36348 ( .A0(n33641), .A1(n33640), .B0(n34696), .C0(n33639), .Y(
        n16393) );
  AOI221XL U36349 ( .A0(n33643), .A1(n16657), .B0(n33642), .B1(n24499), .C0(
        n34763), .Y(n33648) );
  INVXL U36350 ( .A(conv_1[351]), .Y(n33647) );
  OAI211XL U36351 ( .A0(n35441), .A1(n33645), .B0(n32656), .C0(n33644), .Y(
        n33646) );
  OAI211XL U36352 ( .A0(n33648), .A1(n33647), .B0(n34544), .C0(n33646), .Y(
        n16112) );
  AOI221XL U36353 ( .A0(n33651), .A1(n36020), .B0(n33650), .B1(n16656), .C0(
        n33649), .Y(n33657) );
  OAI211XL U36354 ( .A0(n33654), .A1(n33653), .B0(n33778), .C0(n33652), .Y(
        n33655) );
  OAI211XL U36355 ( .A0(n33657), .A1(n33656), .B0(n16652), .C0(n33655), .Y(
        n16063) );
  AOI221XL U36356 ( .A0(n33660), .A1(n36020), .B0(n33659), .B1(n36020), .C0(
        n33658), .Y(n33666) );
  OAI211XL U36357 ( .A0(n33663), .A1(n33662), .B0(n28751), .C0(n33661), .Y(
        n33664) );
  OAI211XL U36358 ( .A0(n33666), .A1(n33665), .B0(n34544), .C0(n33664), .Y(
        n16211) );
  AOI21XL U36359 ( .A0(n34133), .A1(n34132), .B0(n33668), .Y(n33670) );
  NAND2XL U36360 ( .A(conv_2[492]), .B(n33670), .Y(n33669) );
  OAI211XL U36361 ( .A0(conv_2[492]), .A1(n33670), .B0(n16656), .C0(n33669), 
        .Y(n33671) );
  OAI211XL U36362 ( .A0(n34137), .A1(n34131), .B0(n34669), .C0(n33671), .Y(
        n14876) );
  AOI221XL U36363 ( .A0(n33673), .A1(n33712), .B0(n33672), .B1(n16657), .C0(
        n34531), .Y(n33678) );
  INVXL U36364 ( .A(conv_2[383]), .Y(n33677) );
  OAI211XL U36365 ( .A0(n34529), .A1(n33675), .B0(n33982), .C0(n33674), .Y(
        n33676) );
  OAI211XL U36366 ( .A0(n33678), .A1(n33677), .B0(n35859), .C0(n33676), .Y(
        n14950) );
  AOI221XL U36367 ( .A0(n33681), .A1(n33778), .B0(n33680), .B1(n24499), .C0(
        n33679), .Y(n33686) );
  OAI211XL U36368 ( .A0(n35942), .A1(n33683), .B0(n32611), .C0(n33682), .Y(
        n33684) );
  OAI211XL U36369 ( .A0(n33686), .A1(n33685), .B0(n33815), .C0(n33684), .Y(
        n15039) );
  AOI221XL U36370 ( .A0(n33689), .A1(n16656), .B0(n33688), .B1(n36020), .C0(
        n33687), .Y(n33694) );
  OAI211XL U36371 ( .A0(n36045), .A1(n33691), .B0(n33788), .C0(n33690), .Y(
        n33692) );
  OAI211XL U36372 ( .A0(n33694), .A1(n33693), .B0(n34735), .C0(n33692), .Y(
        n14929) );
  NAND3XL U36373 ( .A(n33696), .B(conv_3[402]), .C(n33695), .Y(n34005) );
  NAND3XL U36374 ( .A(n33699), .B(n33698), .C(n33697), .Y(n34004) );
  NAND2XL U36375 ( .A(n34005), .B(n34004), .Y(n33701) );
  NAND2XL U36376 ( .A(conv_3[403]), .B(n33701), .Y(n33700) );
  OAI211XL U36377 ( .A0(conv_3[403]), .A1(n33701), .B0(n33157), .C0(n33700), 
        .Y(n33702) );
  OAI211XL U36378 ( .A0(n33703), .A1(n34003), .B0(n16649), .C0(n33702), .Y(
        n15475) );
  NAND4XL U36379 ( .A(conv_2[506]), .B(conv_2[507]), .C(n36081), .D(n33704), 
        .Y(n34012) );
  NAND2XL U36380 ( .A(n34012), .B(n34011), .Y(n33707) );
  NAND2XL U36381 ( .A(conv_2[508]), .B(n33707), .Y(n33706) );
  OAI211XL U36382 ( .A0(conv_2[508]), .A1(n33707), .B0(n34666), .C0(n33706), 
        .Y(n33708) );
  OAI211XL U36383 ( .A0(n36091), .A1(n34010), .B0(n34669), .C0(n33708), .Y(
        n14865) );
  AOI22XL U36384 ( .A0(n33712), .A1(n33711), .B0(conv_3[132]), .B1(n35572), 
        .Y(n33713) );
  NAND2XL U36385 ( .A(n33713), .B(n35588), .Y(n15656) );
  AOI221XL U36386 ( .A0(n33716), .A1(n33778), .B0(n33715), .B1(n33712), .C0(
        n33714), .Y(n33722) );
  INVXL U36387 ( .A(conv_3[533]), .Y(n33721) );
  OAI211XL U36388 ( .A0(n33719), .A1(n33718), .B0(n33788), .C0(n33717), .Y(
        n33720) );
  OAI211XL U36389 ( .A0(n33722), .A1(n33721), .B0(n35588), .C0(n33720), .Y(
        n15390) );
  AOI221XL U36390 ( .A0(n33724), .A1(n33157), .B0(n33723), .B1(n31735), .C0(
        n33747), .Y(n33729) );
  OAI211XL U36391 ( .A0(n33752), .A1(n33726), .B0(n31735), .C0(n33725), .Y(
        n33727) );
  OAI211XL U36392 ( .A0(n33729), .A1(n33728), .B0(n33468), .C0(n33727), .Y(
        n15506) );
  AOI221XL U36393 ( .A0(n33732), .A1(n24499), .B0(n33731), .B1(n33157), .C0(
        n33730), .Y(n33738) );
  OAI211XL U36394 ( .A0(n33735), .A1(n33734), .B0(n34666), .C0(n33733), .Y(
        n33736) );
  OAI211XL U36395 ( .A0(n33738), .A1(n33737), .B0(n33815), .C0(n33736), .Y(
        n15156) );
  AOI221XL U36396 ( .A0(n33741), .A1(n36020), .B0(n33740), .B1(n31735), .C0(
        n33739), .Y(n33746) );
  INVXL U36397 ( .A(conv_3[96]), .Y(n33745) );
  OAI211XL U36398 ( .A0(n34186), .A1(n33743), .B0(n33778), .C0(n33742), .Y(
        n33744) );
  OAI211XL U36399 ( .A0(n33746), .A1(n33745), .B0(n33468), .C0(n33744), .Y(
        n15682) );
  AOI221XL U36400 ( .A0(n33749), .A1(n16657), .B0(n33748), .B1(n16657), .C0(
        n33747), .Y(n33755) );
  INVXL U36401 ( .A(conv_3[353]), .Y(n33754) );
  OAI211XL U36402 ( .A0(n33752), .A1(n33751), .B0(n33778), .C0(n33750), .Y(
        n33753) );
  OAI211XL U36403 ( .A0(n33755), .A1(n33754), .B0(n16649), .C0(n33753), .Y(
        n15510) );
  AOI221XL U36404 ( .A0(n33758), .A1(n16657), .B0(n33757), .B1(n31735), .C0(
        n33756), .Y(n33764) );
  OAI211XL U36405 ( .A0(n33761), .A1(n33760), .B0(n33788), .C0(n33759), .Y(
        n33762) );
  OAI211XL U36406 ( .A0(n33764), .A1(n33763), .B0(n16649), .C0(n33762), .Y(
        n15448) );
  AOI221XL U36407 ( .A0(n33767), .A1(n24378), .B0(n33766), .B1(n33157), .C0(
        n33765), .Y(n33773) );
  INVXL U36408 ( .A(conv_2[218]), .Y(n33772) );
  OAI211XL U36409 ( .A0(n33770), .A1(n33769), .B0(n34666), .C0(n33768), .Y(
        n33771) );
  OAI211XL U36410 ( .A0(n33773), .A1(n33772), .B0(n35859), .C0(n33771), .Y(
        n15060) );
  AOI221XL U36411 ( .A0(n33776), .A1(n31735), .B0(n33775), .B1(n36020), .C0(
        n33774), .Y(n33783) );
  OAI211XL U36412 ( .A0(n33780), .A1(n33779), .B0(n33778), .C0(n33777), .Y(
        n33781) );
  OAI211XL U36413 ( .A0(n33783), .A1(n33782), .B0(n16649), .C0(n33781), .Y(
        n15441) );
  AOI221XL U36414 ( .A0(n33786), .A1(n33788), .B0(n33785), .B1(n36020), .C0(
        n33784), .Y(n33793) );
  INVXL U36415 ( .A(conv_3[426]), .Y(n33792) );
  OAI211XL U36416 ( .A0(n33790), .A1(n33789), .B0(n33788), .C0(n33787), .Y(
        n33791) );
  OAI211XL U36417 ( .A0(n33793), .A1(n33792), .B0(n16649), .C0(n33791), .Y(
        n15462) );
  AOI221XL U36418 ( .A0(n33795), .A1(n16656), .B0(n33794), .B1(n33712), .C0(
        n35572), .Y(n33800) );
  OAI211XL U36419 ( .A0(n35622), .A1(n33797), .B0(n33778), .C0(n33796), .Y(
        n33798) );
  OAI211XL U36420 ( .A0(n33800), .A1(n33799), .B0(n33468), .C0(n33798), .Y(
        n15658) );
  AOI221XL U36421 ( .A0(n33803), .A1(n16656), .B0(n33802), .B1(n24499), .C0(
        n33801), .Y(n33808) );
  INVXL U36422 ( .A(conv_2[126]), .Y(n33807) );
  OAI211XL U36423 ( .A0(n34344), .A1(n33805), .B0(n33778), .C0(n33804), .Y(
        n33806) );
  OAI211XL U36424 ( .A0(n33808), .A1(n33807), .B0(n33815), .C0(n33806), .Y(
        n15122) );
  AOI221XL U36425 ( .A0(n33811), .A1(n33778), .B0(n33810), .B1(n36020), .C0(
        n33809), .Y(n33817) );
  OAI211XL U36426 ( .A0(n35876), .A1(n33813), .B0(n33788), .C0(n33812), .Y(
        n33814) );
  OAI211XL U36427 ( .A0(n33817), .A1(n33816), .B0(n33815), .C0(n33814), .Y(
        n15148) );
  AOI221XL U36428 ( .A0(n33820), .A1(n28751), .B0(n33819), .B1(n33788), .C0(
        n33818), .Y(n33827) );
  INVXL U36429 ( .A(conv_3[57]), .Y(n33826) );
  OAI211XL U36430 ( .A0(n33824), .A1(n33823), .B0(n33822), .C0(n33821), .Y(
        n33825) );
  OAI211XL U36431 ( .A0(n33827), .A1(n33826), .B0(n33468), .C0(n33825), .Y(
        n15706) );
  AOI221XL U36432 ( .A0(n33830), .A1(n33788), .B0(n33829), .B1(n36020), .C0(
        n33828), .Y(n33836) );
  OAI211XL U36433 ( .A0(n33833), .A1(n33832), .B0(n16657), .C0(n33831), .Y(
        n33834) );
  OAI211XL U36434 ( .A0(n33836), .A1(n33835), .B0(n33468), .C0(n33834), .Y(
        n15498) );
  AOI221XL U36435 ( .A0(n33839), .A1(n34028), .B0(n33838), .B1(n24499), .C0(
        n33837), .Y(n33845) );
  INVXL U36436 ( .A(conv_3[322]), .Y(n33844) );
  OAI211XL U36437 ( .A0(n33842), .A1(n33841), .B0(n30090), .C0(n33840), .Y(
        n33843) );
  OAI211XL U36438 ( .A0(n33845), .A1(n33844), .B0(n16649), .C0(n33843), .Y(
        n15531) );
  AOI22XL U36439 ( .A0(conv_1[238]), .A1(n33848), .B0(n33847), .B1(n33846), 
        .Y(n33850) );
  NAND2XL U36440 ( .A(conv_1[239]), .B(n33850), .Y(n33849) );
  OAI211XL U36441 ( .A0(conv_1[239]), .A1(n33850), .B0(n33778), .C0(n33849), 
        .Y(n33851) );
  OAI211XL U36442 ( .A0(n33853), .A1(n33852), .B0(n34281), .C0(n33851), .Y(
        n16224) );
  INVXL U36443 ( .A(conv_3[507]), .Y(n33920) );
  NAND2XL U36444 ( .A(n33855), .B(n33854), .Y(n33856) );
  AOI32XL U36445 ( .A0(conv_3[506]), .A1(n33919), .A2(n33917), .B0(n35838), 
        .B1(n33919), .Y(n33858) );
  NAND2XL U36446 ( .A(n33920), .B(n33858), .Y(n33857) );
  OAI211XL U36447 ( .A0(n33920), .A1(n33858), .B0(n33982), .C0(n33857), .Y(
        n33859) );
  OAI211XL U36448 ( .A0(n35841), .A1(n33920), .B0(n16649), .C0(n33859), .Y(
        n15406) );
  OAI21XL U36449 ( .A0(n33860), .A1(n16654), .B0(n34263), .Y(n33861) );
  AOI32XL U36450 ( .A0(n34465), .A1(n33861), .A2(n34769), .B0(conv_1[315]), 
        .B1(n33861), .Y(n33862) );
  NAND2XL U36451 ( .A(n34773), .B(n33862), .Y(n16148) );
  OAI2BB1XL U36452 ( .A0N(n36020), .A1N(n33864), .B0(n33863), .Y(n33865) );
  AOI32XL U36453 ( .A0(n33867), .A1(n33866), .A2(n34769), .B0(conv_1[300]), 
        .B1(n33865), .Y(n33868) );
  NAND2XL U36454 ( .A(n33868), .B(n34773), .Y(n16163) );
  OAI21XL U36455 ( .A0(n33869), .A1(n16655), .B0(n35395), .Y(n33870) );
  AOI32XL U36456 ( .A0(n34476), .A1(n33871), .A2(n34769), .B0(conv_1[210]), 
        .B1(n33870), .Y(n33872) );
  NAND2XL U36457 ( .A(n33872), .B(n34773), .Y(n16253) );
  OAI21XL U36458 ( .A0(n33873), .A1(n16654), .B0(n35408), .Y(n33874) );
  AOI32XL U36459 ( .A0(n34461), .A1(n33875), .A2(n34769), .B0(conv_1[225]), 
        .B1(n33874), .Y(n33876) );
  NAND2XL U36460 ( .A(n33876), .B(n34773), .Y(n16238) );
  NAND4XL U36461 ( .A(conv_3[236]), .B(conv_3[237]), .C(n33878), .D(n33877), 
        .Y(n33900) );
  NAND3XL U36462 ( .A(n35673), .B(n33880), .C(n33879), .Y(n33899) );
  NAND2XL U36463 ( .A(n33900), .B(n33899), .Y(n33882) );
  OAI21XL U36464 ( .A0(n16654), .A1(n33882), .B0(n35676), .Y(n33881) );
  NAND2XL U36465 ( .A(n33883), .B(n35588), .Y(n15585) );
  AOI32XL U36466 ( .A0(conv_1[341]), .A1(n33885), .A2(n33884), .B0(n35434), 
        .B1(n33885), .Y(n33887) );
  AOI211XL U36467 ( .A0(n33889), .A1(n33887), .B0(n16654), .C0(n33886), .Y(
        n33888) );
  AOI2BB1XL U36468 ( .A0N(n33889), .A1N(n35437), .B0(n33888), .Y(n33890) );
  NAND2XL U36469 ( .A(n33890), .B(n34544), .Y(n16121) );
  NAND2XL U36470 ( .A(n33892), .B(n33891), .Y(n33894) );
  AOI211XL U36471 ( .A0(n33896), .A1(n33894), .B0(n36009), .C0(n33893), .Y(
        n33895) );
  NAND2XL U36472 ( .A(n33897), .B(n34735), .Y(n14893) );
  AOI22XL U36473 ( .A0(conv_3[238]), .A1(n33900), .B0(n33899), .B1(n33898), 
        .Y(n33902) );
  NAND2XL U36474 ( .A(conv_3[239]), .B(n33902), .Y(n33901) );
  OAI211XL U36475 ( .A0(conv_3[239]), .A1(n33902), .B0(n33778), .C0(n33901), 
        .Y(n33903) );
  OAI211XL U36476 ( .A0(n34789), .A1(n33904), .B0(n35588), .C0(n33903), .Y(
        n15584) );
  OAI211XL U36477 ( .A0(conv_3[269]), .A1(n33909), .B0(n33788), .C0(n33908), 
        .Y(n33910) );
  INVXL U36478 ( .A(conv_3[30]), .Y(n33915) );
  AOI32XL U36479 ( .A0(n33913), .A1(n35594), .A2(n33990), .B0(n16654), .B1(
        n35594), .Y(n33914) );
  AOI32XL U36480 ( .A0(n34742), .A1(n33915), .A2(n33990), .B0(conv_3[30]), 
        .B1(n33914), .Y(n33916) );
  NAND2XL U36481 ( .A(n33916), .B(n34755), .Y(n15921) );
  INVXL U36482 ( .A(conv_3[508]), .Y(n34513) );
  NAND4XL U36483 ( .A(conv_3[506]), .B(conv_3[507]), .C(n33918), .D(n33917), 
        .Y(n34515) );
  NAND3XL U36484 ( .A(n35838), .B(n33920), .C(n33919), .Y(n34514) );
  NAND2XL U36485 ( .A(n34515), .B(n34514), .Y(n33922) );
  NAND2XL U36486 ( .A(conv_3[508]), .B(n33922), .Y(n33921) );
  OAI211XL U36487 ( .A0(conv_3[508]), .A1(n33922), .B0(n27932), .C0(n33921), 
        .Y(n33923) );
  OAI211XL U36488 ( .A0(n35841), .A1(n34513), .B0(n16649), .C0(n33923), .Y(
        n15405) );
  NAND2XL U36489 ( .A(n33925), .B(n33924), .Y(n33927) );
  NAND2XL U36490 ( .A(n33927), .B(n33926), .Y(n33929) );
  AOI211XL U36491 ( .A0(n33931), .A1(n33929), .B0(n16658), .C0(n33928), .Y(
        n33930) );
  AOI2BB1XL U36492 ( .A0N(n33931), .A1N(n36010), .B0(n33930), .Y(n33932) );
  NAND2XL U36493 ( .A(n33932), .B(n35859), .Y(n14973) );
  AOI32XL U36494 ( .A0(conv_2[326]), .A1(n33934), .A2(n33933), .B0(n35982), 
        .B1(n33934), .Y(n33936) );
  AOI211XL U36495 ( .A0(n33938), .A1(n33936), .B0(n36009), .C0(n33935), .Y(
        n33937) );
  NAND2XL U36496 ( .A(n33939), .B(n35859), .Y(n14986) );
  NAND2XL U36497 ( .A(n33940), .B(n33946), .Y(n33942) );
  AOI211XL U36498 ( .A0(n33944), .A1(n33942), .B0(n16655), .C0(n33941), .Y(
        n33943) );
  NAND2XL U36499 ( .A(n33945), .B(n35859), .Y(n15097) );
  AOI32XL U36500 ( .A0(conv_2[161]), .A1(n33947), .A2(n33946), .B0(n34626), 
        .B1(n33947), .Y(n33949) );
  AOI211XL U36501 ( .A0(n33951), .A1(n33949), .B0(n16655), .C0(n33948), .Y(
        n33950) );
  NAND2XL U36502 ( .A(n33952), .B(n35859), .Y(n15096) );
  AOI32XL U36503 ( .A0(conv_2[401]), .A1(n33953), .A2(n36033), .B0(n34634), 
        .B1(n36034), .Y(n33955) );
  AOI211XL U36504 ( .A0(n33957), .A1(n33955), .B0(n16655), .C0(n33954), .Y(
        n33956) );
  AOI2BB1XL U36505 ( .A0N(n33957), .A1N(n36031), .B0(n33956), .Y(n33958) );
  NAND2XL U36506 ( .A(n33958), .B(n35859), .Y(n14936) );
  OAI21XL U36507 ( .A0(n35831), .A1(n33960), .B0(n33959), .Y(n33962) );
  AOI211XL U36508 ( .A0(n33964), .A1(n33962), .B0(n16655), .C0(n33961), .Y(
        n33963) );
  AOI2BB1XL U36509 ( .A0N(n33964), .A1N(n35826), .B0(n33963), .Y(n33965) );
  NAND2XL U36510 ( .A(n33965), .B(n35588), .Y(n15420) );
  NAND2BXL U36511 ( .AN(n33967), .B(n33966), .Y(n33969) );
  AOI211XL U36512 ( .A0(n33971), .A1(n33969), .B0(n16655), .C0(n33968), .Y(
        n33970) );
  AOI2BB1XL U36513 ( .A0N(n33971), .A1N(n34737), .B0(n33970), .Y(n33972) );
  NAND2XL U36514 ( .A(n33972), .B(n35588), .Y(n15647) );
  INVXL U36515 ( .A(conv_2[178]), .Y(n34592) );
  ADDFX1 U36516 ( .A(conv_2[176]), .B(n29831), .CI(n33973), .CO(n34585), .S(
        n30898) );
  NAND3XL U36517 ( .A(conv_2[177]), .B(n34585), .C(n33974), .Y(n34594) );
  NAND2XL U36518 ( .A(n34594), .B(n34593), .Y(n33976) );
  NAND2XL U36519 ( .A(conv_2[178]), .B(n33976), .Y(n33975) );
  OAI211XL U36520 ( .A0(conv_2[178]), .A1(n33976), .B0(n16657), .C0(n33975), 
        .Y(n33977) );
  OAI211XL U36521 ( .A0(n34589), .A1(n34592), .B0(n35859), .C0(n33977), .Y(
        n15085) );
  ADDFX1 U36522 ( .A(conv_2[312]), .B(n33979), .CI(n33978), .CO(n33980), .S(
        n28629) );
  NOR2X1 U36523 ( .A(n33980), .B(n35970), .Y(n34024) );
  NOR2X1 U36524 ( .A(conv_2[313]), .B(n34024), .Y(n34023) );
  AOI21XL U36525 ( .A0(conv_2[313]), .A1(n34022), .B0(n34023), .Y(n33983) );
  NAND2XL U36526 ( .A(conv_2[314]), .B(n33983), .Y(n33981) );
  OAI211XL U36527 ( .A0(conv_2[314]), .A1(n33983), .B0(n33982), .C0(n33981), 
        .Y(n33984) );
  OAI211XL U36528 ( .A0(n33442), .A1(n33985), .B0(n33815), .C0(n33984), .Y(
        n14994) );
  AOI221XL U36529 ( .A0(n33988), .A1(n34028), .B0(n33987), .B1(n33778), .C0(
        n33986), .Y(n33992) );
  AOI21XL U36530 ( .A0(n34581), .A1(n33990), .B0(conv_2[30]), .Y(n33991) );
  OAI21XL U36531 ( .A0(n33992), .A1(n33991), .B0(n34583), .Y(n15381) );
  AOI221XL U36532 ( .A0(n33994), .A1(n32611), .B0(n33993), .B1(n35336), .C0(
        n35952), .Y(n33996) );
  AOI21XL U36533 ( .A0(n34581), .A1(n34711), .B0(conv_2[270]), .Y(n33995) );
  OAI21XL U36534 ( .A0(n33996), .A1(n33995), .B0(n34583), .Y(n15365) );
  NAND2XL U36535 ( .A(n33998), .B(n33997), .Y(n34000) );
  OAI21XL U36536 ( .A0(n35419), .A1(n34000), .B0(n35447), .Y(n33999) );
  AOI32XL U36537 ( .A0(n36020), .A1(n34001), .A2(n34000), .B0(conv_1[358]), 
        .B1(n33999), .Y(n34002) );
  NAND2XL U36538 ( .A(n34002), .B(n34281), .Y(n16105) );
  AOI22XL U36539 ( .A0(conv_3[403]), .A1(n34005), .B0(n34004), .B1(n34003), 
        .Y(n34007) );
  NAND2XL U36540 ( .A(conv_3[404]), .B(n34007), .Y(n34006) );
  OAI211XL U36541 ( .A0(conv_3[404]), .A1(n34007), .B0(n33778), .C0(n34006), 
        .Y(n34008) );
  OAI211XL U36542 ( .A0(n34520), .A1(n34009), .B0(n33468), .C0(n34008), .Y(
        n15474) );
  AOI22XL U36543 ( .A0(conv_2[508]), .A1(n34012), .B0(n34011), .B1(n34010), 
        .Y(n34014) );
  NAND2XL U36544 ( .A(conv_2[509]), .B(n34014), .Y(n34013) );
  OAI211XL U36545 ( .A0(conv_2[509]), .A1(n34014), .B0(n32611), .C0(n34013), 
        .Y(n34015) );
  OAI211XL U36546 ( .A0(n34676), .A1(n34016), .B0(n34669), .C0(n34015), .Y(
        n14864) );
  INVXL U36547 ( .A(conv_1[510]), .Y(n34020) );
  AOI32XL U36548 ( .A0(n34017), .A1(n35547), .A2(n34019), .B0(n34389), .B1(
        n35547), .Y(n34018) );
  AOI32XL U36549 ( .A0(n34769), .A1(n34020), .A2(n34019), .B0(conv_1[510]), 
        .B1(n34018), .Y(n34021) );
  NAND2XL U36550 ( .A(n34021), .B(n34773), .Y(n15953) );
  INVXL U36551 ( .A(n34022), .Y(n34025) );
  AOI22XL U36552 ( .A0(n34028), .A1(n34027), .B0(conv_2[313]), .B1(n34026), 
        .Y(n34029) );
  NAND2XL U36553 ( .A(n34029), .B(n35859), .Y(n14995) );
  OAI21XL U36554 ( .A0(n35419), .A1(n34033), .B0(n35736), .Y(n34032) );
  NAND2XL U36555 ( .A(n34035), .B(n16649), .Y(n15535) );
  OAI21XL U36556 ( .A0(n35419), .A1(n34039), .B0(n36047), .Y(n34038) );
  NAND2XL U36557 ( .A(n34041), .B(n34735), .Y(n14925) );
  INVXL U36558 ( .A(conv_1[158]), .Y(n34049) );
  NAND2XL U36559 ( .A(n34044), .B(n34043), .Y(n34042) );
  OAI21XL U36560 ( .A0(n34044), .A1(n34043), .B0(n34042), .Y(n34046) );
  AOI211XL U36561 ( .A0(n34049), .A1(n34046), .B0(n16655), .C0(n34045), .Y(
        n34047) );
  NAND2XL U36562 ( .A(n34050), .B(n34682), .Y(n16305) );
  OAI21XL U36563 ( .A0(n34053), .A1(n34052), .B0(n34051), .Y(n34055) );
  AOI211XL U36564 ( .A0(n34058), .A1(n34055), .B0(n36009), .C0(n34054), .Y(
        n34056) );
  NAND2XL U36565 ( .A(n34059), .B(n34281), .Y(n16381) );
  AOI32XL U36566 ( .A0(conv_1[206]), .A1(n34060), .A2(n35386), .B0(n35379), 
        .B1(n35387), .Y(n34062) );
  AOI211XL U36567 ( .A0(n34064), .A1(n34062), .B0(n16655), .C0(n34061), .Y(
        n34063) );
  NAND2XL U36568 ( .A(n34065), .B(n34544), .Y(n16256) );
  OAI21XL U36569 ( .A0(n35419), .A1(n34069), .B0(n35743), .Y(n34068) );
  NAND2XL U36570 ( .A(n34071), .B(n16649), .Y(n15525) );
  INVXL U36571 ( .A(conv_3[424]), .Y(n34076) );
  OAI21XL U36572 ( .A0(n34075), .A1(n16655), .B0(n35778), .Y(n34074) );
  NAND2XL U36573 ( .A(n34077), .B(n34097), .Y(n15751) );
  NAND2XL U36574 ( .A(n34079), .B(n34078), .Y(n34082) );
  OAI21XL U36575 ( .A0(n16654), .A1(n34082), .B0(n34080), .Y(n34081) );
  NAND2XL U36576 ( .A(n34084), .B(n34544), .Y(n16195) );
  AOI32XL U36577 ( .A0(conv_1[191]), .A1(n34086), .A2(n34085), .B0(n35365), 
        .B1(n34086), .Y(n34088) );
  AOI211XL U36578 ( .A0(n34090), .A1(n34088), .B0(n35419), .C0(n34087), .Y(
        n34089) );
  NAND2XL U36579 ( .A(n34091), .B(n34689), .Y(n16271) );
  INVXL U36580 ( .A(conv_3[499]), .Y(n34096) );
  OAI21XL U36581 ( .A0(n34095), .A1(n35419), .B0(n35841), .Y(n34094) );
  NAND2XL U36582 ( .A(n34098), .B(n34097), .Y(n15746) );
  NAND2XL U36583 ( .A(n34100), .B(n34099), .Y(n34102) );
  AOI211XL U36584 ( .A0(n34104), .A1(n34102), .B0(n16654), .C0(n34101), .Y(
        n34103) );
  NAND2XL U36585 ( .A(n34106), .B(n34105), .Y(n15242) );
  NAND2XL U36586 ( .A(n34108), .B(n34107), .Y(n34110) );
  AOI211XL U36587 ( .A0(n34112), .A1(n34110), .B0(n34389), .C0(n34109), .Y(
        n34111) );
  NAND2XL U36588 ( .A(n34113), .B(n35574), .Y(n15811) );
  INVXL U36589 ( .A(conv_2[195]), .Y(n34116) );
  OAI21XL U36590 ( .A0(n16654), .A1(n34115), .B0(n35931), .Y(n34114) );
  AOI32XL U36591 ( .A0(n36020), .A1(n34116), .A2(n34115), .B0(conv_2[195]), 
        .B1(n34114), .Y(n34117) );
  NAND2XL U36592 ( .A(n34117), .B(n34583), .Y(n15370) );
  OAI21XL U36593 ( .A0(n35419), .A1(n34121), .B0(n35368), .Y(n34120) );
  NAND2XL U36594 ( .A(n34123), .B(n34281), .Y(n16270) );
  OAI21XL U36595 ( .A0(n34127), .A1(n16654), .B0(n34491), .Y(n34126) );
  AOI32XL U36596 ( .A0(n36020), .A1(n34128), .A2(n34127), .B0(conv_2[125]), 
        .B1(n34126), .Y(n34129) );
  NAND2XL U36597 ( .A(n34129), .B(n34735), .Y(n15123) );
  NAND3XL U36598 ( .A(conv_2[492]), .B(n34133), .C(n34130), .Y(n34664) );
  NAND2XL U36599 ( .A(n34664), .B(n34663), .Y(n34135) );
  NAND2XL U36600 ( .A(conv_2[493]), .B(n34135), .Y(n34134) );
  OAI211XL U36601 ( .A0(conv_2[493]), .A1(n34135), .B0(n34666), .C0(n34134), 
        .Y(n34136) );
  OAI211XL U36602 ( .A0(n34137), .A1(n34662), .B0(n34669), .C0(n34136), .Y(
        n14875) );
  OAI21XL U36603 ( .A0(n16655), .A1(n34141), .B0(n34168), .Y(n34140) );
  NAND2XL U36604 ( .A(n34143), .B(n16649), .Y(n15485) );
  NAND2XL U36605 ( .A(n34145), .B(n34144), .Y(n34147) );
  OAI21XL U36606 ( .A0(n16654), .A1(n34147), .B0(n35945), .Y(n34146) );
  NAND2XL U36607 ( .A(n34149), .B(n35859), .Y(n15035) );
  OAI21XL U36608 ( .A0(n34153), .A1(n36009), .B0(n35610), .Y(n34152) );
  AOI32XL U36609 ( .A0(n33982), .A1(n34154), .A2(n34153), .B0(conv_3[80]), 
        .B1(n34152), .Y(n34155) );
  NAND2XL U36610 ( .A(n34155), .B(n16649), .Y(n15693) );
  NAND2XL U36611 ( .A(n34157), .B(n34156), .Y(n34159) );
  OAI21XL U36612 ( .A0(n16655), .A1(n34159), .B0(n34392), .Y(n34158) );
  NAND2XL U36613 ( .A(n34161), .B(n16649), .Y(n15705) );
  OAI21XL U36614 ( .A0(n34164), .A1(n34163), .B0(n34162), .Y(n34166) );
  AOI211XL U36615 ( .A0(n34169), .A1(n34166), .B0(n16654), .C0(n34165), .Y(
        n34167) );
  NAND2XL U36616 ( .A(n34170), .B(n16649), .Y(n15486) );
  OAI21XL U36617 ( .A0(n34173), .A1(n34172), .B0(n34171), .Y(n34175) );
  AOI211XL U36618 ( .A0(n34178), .A1(n34175), .B0(n16658), .C0(n34174), .Y(
        n34176) );
  NAND2XL U36619 ( .A(n34179), .B(n34735), .Y(n14888) );
  NAND2XL U36620 ( .A(n34180), .B(n34187), .Y(n34182) );
  AOI211XL U36621 ( .A0(n34184), .A1(n34182), .B0(n34389), .C0(n34181), .Y(
        n34183) );
  NAND2XL U36622 ( .A(n34185), .B(n16649), .Y(n15677) );
  AOI32XL U36623 ( .A0(conv_3[101]), .A1(n34188), .A2(n34187), .B0(n34186), 
        .B1(n34188), .Y(n34190) );
  AOI211XL U36624 ( .A0(n34192), .A1(n34190), .B0(n34389), .C0(n34189), .Y(
        n34191) );
  NAND2XL U36625 ( .A(n34193), .B(n16649), .Y(n15676) );
  OAI21XL U36626 ( .A0(n34196), .A1(n34195), .B0(n34194), .Y(n34198) );
  AOI211XL U36627 ( .A0(n34201), .A1(n34198), .B0(n34389), .C0(n34197), .Y(
        n34199) );
  NAND2XL U36628 ( .A(n34202), .B(n16649), .Y(n15666) );
  INVXL U36629 ( .A(conv_2[432]), .Y(n34207) );
  OAI21XL U36630 ( .A0(conv_2[431]), .A1(n34210), .B0(n34211), .Y(n34203) );
  AOI32XL U36631 ( .A0(conv_2[431]), .A1(n34203), .A2(n34210), .B0(n34211), 
        .B1(n34203), .Y(n34205) );
  AOI211XL U36632 ( .A0(n34207), .A1(n34205), .B0(n35419), .C0(n34204), .Y(
        n34206) );
  NAND2XL U36633 ( .A(n34208), .B(n34735), .Y(n14916) );
  INVXL U36634 ( .A(conv_2[431]), .Y(n34215) );
  NAND2XL U36635 ( .A(n34211), .B(n34210), .Y(n34209) );
  OAI21XL U36636 ( .A0(n34211), .A1(n34210), .B0(n34209), .Y(n34213) );
  AOI211XL U36637 ( .A0(n34215), .A1(n34213), .B0(n16654), .C0(n34212), .Y(
        n34214) );
  NAND2XL U36638 ( .A(n34216), .B(n34735), .Y(n14917) );
  NAND2XL U36639 ( .A(n34218), .B(n34217), .Y(n34220) );
  OAI21XL U36640 ( .A0(n35419), .A1(n34220), .B0(n36003), .Y(n34219) );
  AOI32XL U36641 ( .A0(n33822), .A1(n34221), .A2(n34220), .B0(conv_2[343]), 
        .B1(n34219), .Y(n34222) );
  NAND2XL U36642 ( .A(n34222), .B(n35859), .Y(n14975) );
  AOI32XL U36643 ( .A0(n34223), .A1(n35792), .A2(n34224), .B0(n16654), .B1(
        n35792), .Y(n34225) );
  AOI32XL U36644 ( .A0(n34742), .A1(n34225), .A2(n34224), .B0(conv_3[435]), 
        .B1(n34225), .Y(n34226) );
  NAND2XL U36645 ( .A(n34755), .B(n34226), .Y(n15894) );
  AOI32XL U36646 ( .A0(n34228), .A1(n34227), .A2(n34229), .B0(n35419), .B1(
        n34227), .Y(n34230) );
  AOI32XL U36647 ( .A0(n34742), .A1(n34230), .A2(n34229), .B0(conv_3[405]), 
        .B1(n34230), .Y(n34231) );
  NAND2XL U36648 ( .A(n34755), .B(n34231), .Y(n15896) );
  NAND2BXL U36649 ( .AN(n34233), .B(n34232), .Y(n34235) );
  AOI211XL U36650 ( .A0(n34237), .A1(n34235), .B0(n34389), .C0(n34234), .Y(
        n34236) );
  NAND2XL U36651 ( .A(n34238), .B(n35847), .Y(n15314) );
  OAI21XL U36652 ( .A0(n34242), .A1(n34389), .B0(n35902), .Y(n34241) );
  AOI32XL U36653 ( .A0(n34028), .A1(n34243), .A2(n34242), .B0(conv_2[140]), 
        .B1(n34241), .Y(n34244) );
  NAND2XL U36654 ( .A(n34244), .B(n35859), .Y(n15113) );
  OAI21XL U36655 ( .A0(n34248), .A1(n16654), .B0(n35706), .Y(n34247) );
  NAND2XL U36656 ( .A(n34250), .B(n35588), .Y(n15583) );
  INVXL U36657 ( .A(conv_1[327]), .Y(n34255) );
  OAI21XL U36658 ( .A0(conv_1[326]), .A1(n34258), .B0(n34259), .Y(n34251) );
  AOI32XL U36659 ( .A0(conv_1[326]), .A1(n34251), .A2(n34258), .B0(n34259), 
        .B1(n34251), .Y(n34253) );
  AOI211XL U36660 ( .A0(n34255), .A1(n34253), .B0(n36042), .C0(n34252), .Y(
        n34254) );
  NAND2XL U36661 ( .A(n34256), .B(n34544), .Y(n16136) );
  INVXL U36662 ( .A(conv_1[326]), .Y(n34264) );
  NAND2XL U36663 ( .A(n34259), .B(n34258), .Y(n34257) );
  OAI21XL U36664 ( .A0(n34259), .A1(n34258), .B0(n34257), .Y(n34261) );
  AOI211XL U36665 ( .A0(n34264), .A1(n34261), .B0(n36001), .C0(n34260), .Y(
        n34262) );
  NAND2XL U36666 ( .A(n34265), .B(n34682), .Y(n16137) );
  NAND2XL U36667 ( .A(n34267), .B(n34266), .Y(n34269) );
  AOI211XL U36668 ( .A0(n34272), .A1(n34269), .B0(n36009), .C0(n34268), .Y(
        n34270) );
  NAND2XL U36669 ( .A(n34273), .B(n34682), .Y(n16317) );
  AOI32XL U36670 ( .A0(conv_1[236]), .A1(n34276), .A2(n34275), .B0(n35404), 
        .B1(n34274), .Y(n34278) );
  AOI211XL U36671 ( .A0(n34280), .A1(n34278), .B0(n36001), .C0(n34277), .Y(
        n34279) );
  NAND2XL U36672 ( .A(n34282), .B(n34281), .Y(n16226) );
  NAND2XL U36673 ( .A(n34283), .B(n34306), .Y(n34285) );
  AOI211XL U36674 ( .A0(n34287), .A1(n34285), .B0(n36001), .C0(n34284), .Y(
        n34286) );
  NAND2XL U36675 ( .A(n34288), .B(n34696), .Y(n16092) );
  INVXL U36676 ( .A(conv_1[128]), .Y(n34297) );
  OAI21XL U36677 ( .A0(conv_1[127]), .A1(n34289), .B0(n34292), .Y(n34290) );
  OAI21XL U36678 ( .A0(n34292), .A1(n34291), .B0(n34290), .Y(n34294) );
  AOI211XL U36679 ( .A0(n34297), .A1(n34294), .B0(n36042), .C0(n34293), .Y(
        n34295) );
  NAND2XL U36680 ( .A(n34298), .B(n34696), .Y(n16335) );
  OAI21XL U36681 ( .A0(n35392), .A1(n34300), .B0(n34299), .Y(n34302) );
  AOI211XL U36682 ( .A0(n34304), .A1(n34302), .B0(n35419), .C0(n34301), .Y(
        n34303) );
  NAND2XL U36683 ( .A(n34305), .B(n34544), .Y(n16241) );
  AOI32XL U36684 ( .A0(conv_1[371]), .A1(n34307), .A2(n34306), .B0(n35455), 
        .B1(n34307), .Y(n34309) );
  AOI211XL U36685 ( .A0(n34311), .A1(n34309), .B0(n36009), .C0(n34308), .Y(
        n34310) );
  NAND2XL U36686 ( .A(n34312), .B(n34696), .Y(n16091) );
  NAND2XL U36687 ( .A(n34313), .B(n34320), .Y(n34315) );
  AOI211XL U36688 ( .A0(n34317), .A1(n34315), .B0(n36001), .C0(n34314), .Y(
        n34316) );
  NAND2XL U36689 ( .A(n34318), .B(n34689), .Y(n16167) );
  AOI32XL U36690 ( .A0(conv_1[296]), .A1(n34321), .A2(n34320), .B0(n34319), 
        .B1(n34321), .Y(n34323) );
  AOI211XL U36691 ( .A0(n34326), .A1(n34323), .B0(n36001), .C0(n34322), .Y(
        n34324) );
  NAND2XL U36692 ( .A(n34327), .B(n34689), .Y(n16166) );
  NAND2BXL U36693 ( .AN(n34329), .B(n34328), .Y(n34331) );
  AOI211XL U36694 ( .A0(n34333), .A1(n34331), .B0(n36042), .C0(n34330), .Y(
        n34332) );
  NAND2XL U36695 ( .A(n34334), .B(n34544), .Y(n16217) );
  NAND2BXL U36696 ( .AN(n34336), .B(n34335), .Y(n34338) );
  AOI211XL U36697 ( .A0(n34340), .A1(n34338), .B0(n16654), .C0(n34337), .Y(
        n34339) );
  AOI2BB1XL U36698 ( .A0N(n34340), .A1N(n35466), .B0(n34339), .Y(n34341) );
  NAND2XL U36699 ( .A(n16652), .B(n34341), .Y(n16079) );
  INVXL U36700 ( .A(conv_2[129]), .Y(n34348) );
  NAND2XL U36701 ( .A(n34344), .B(n34343), .Y(n34342) );
  OAI21XL U36702 ( .A0(n34344), .A1(n34343), .B0(n34342), .Y(n34346) );
  AOI211XL U36703 ( .A0(n34348), .A1(n34346), .B0(n34389), .C0(n34345), .Y(
        n34347) );
  NAND2XL U36704 ( .A(n34349), .B(n35859), .Y(n15119) );
  NAND2BXL U36705 ( .AN(n34351), .B(n34350), .Y(n34353) );
  AOI211XL U36706 ( .A0(n34355), .A1(n34353), .B0(n34389), .C0(n34352), .Y(
        n34354) );
  NAND2XL U36707 ( .A(n34356), .B(n35859), .Y(n15117) );
  NAND2XL U36708 ( .A(n34358), .B(n34357), .Y(n34360) );
  AOI211XL U36709 ( .A0(n34362), .A1(n34360), .B0(n34389), .C0(n34359), .Y(
        n34361) );
  NAND2XL U36710 ( .A(n34363), .B(n35859), .Y(n15107) );
  AOI32XL U36711 ( .A0(conv_2[116]), .A1(n34364), .A2(n34642), .B0(n35891), 
        .B1(n34364), .Y(n34366) );
  AOI211XL U36712 ( .A0(n34368), .A1(n34366), .B0(n34389), .C0(n34365), .Y(
        n34367) );
  NAND2XL U36713 ( .A(n34369), .B(n35859), .Y(n15126) );
  NAND2XL U36714 ( .A(n34371), .B(n34370), .Y(n34373) );
  AOI211XL U36715 ( .A0(n34375), .A1(n34373), .B0(n34389), .C0(n34372), .Y(
        n34374) );
  NAND2XL U36716 ( .A(n34376), .B(n35588), .Y(n15713) );
  INVXL U36717 ( .A(conv_3[11]), .Y(n34384) );
  NAND2XL U36718 ( .A(n34379), .B(n34378), .Y(n34377) );
  OAI21XL U36719 ( .A0(n34379), .A1(n34378), .B0(n34377), .Y(n34381) );
  AOI211XL U36720 ( .A0(n34384), .A1(n34381), .B0(n34389), .C0(n34380), .Y(
        n34382) );
  NAND2XL U36721 ( .A(n34385), .B(n35588), .Y(n15737) );
  NAND2XL U36722 ( .A(n34387), .B(n34386), .Y(n34390) );
  AOI211XL U36723 ( .A0(n34393), .A1(n34390), .B0(n34389), .C0(n34388), .Y(
        n34391) );
  NAND2XL U36724 ( .A(n34394), .B(n35588), .Y(n15710) );
  NAND2XL U36725 ( .A(n34396), .B(n34395), .Y(n34398) );
  AOI211XL U36726 ( .A0(n34400), .A1(n34398), .B0(n16654), .C0(n34397), .Y(
        n34399) );
  NAND2XL U36727 ( .A(n34401), .B(n35588), .Y(n15653) );
  NAND2XL U36728 ( .A(n34403), .B(n34402), .Y(n34405) );
  AOI211XL U36729 ( .A0(n34407), .A1(n34405), .B0(n36042), .C0(n34404), .Y(
        n34406) );
  NAND2XL U36730 ( .A(n34409), .B(n34408), .Y(n15232) );
  NAND2XL U36731 ( .A(n34411), .B(n34410), .Y(n34413) );
  OAI21XL U36732 ( .A0(n16654), .A1(n34413), .B0(n35576), .Y(n34412) );
  NAND2XL U36733 ( .A(n34415), .B(n35588), .Y(n15725) );
  OAI2BB1XL U36734 ( .A0N(n36020), .A1N(n34416), .B0(n36010), .Y(n34417) );
  AOI32XL U36735 ( .A0(n34581), .A1(n34418), .A2(n34762), .B0(conv_2[345]), 
        .B1(n34417), .Y(n34419) );
  NAND2XL U36736 ( .A(n34419), .B(n34583), .Y(n15360) );
  INVXL U36737 ( .A(conv_2[255]), .Y(n34423) );
  AOI32XL U36738 ( .A0(n34420), .A1(n34601), .A2(n34422), .B0(n34389), .B1(
        n34601), .Y(n34421) );
  AOI32XL U36739 ( .A0(n34581), .A1(n34423), .A2(n34422), .B0(conv_2[255]), 
        .B1(n34421), .Y(n34424) );
  NAND2XL U36740 ( .A(n34424), .B(n34583), .Y(n15366) );
  INVXL U36741 ( .A(conv_2[135]), .Y(n34429) );
  OAI21XL U36742 ( .A0(n34427), .A1(n34389), .B0(n35902), .Y(n34428) );
  AOI32XL U36743 ( .A0(n34581), .A1(n34429), .A2(n34740), .B0(conv_2[135]), 
        .B1(n34428), .Y(n34430) );
  NAND2XL U36744 ( .A(n34430), .B(n34583), .Y(n15374) );
  OAI21XL U36745 ( .A0(n34431), .A1(n36042), .B0(n34589), .Y(n34432) );
  AOI32XL U36746 ( .A0(n34581), .A1(n34434), .A2(n34433), .B0(conv_2[165]), 
        .B1(n34432), .Y(n34435) );
  NAND2XL U36747 ( .A(n34435), .B(n34583), .Y(n15372) );
  AOI32XL U36748 ( .A0(n34436), .A1(n35879), .A2(n34438), .B0(n36001), .B1(
        n35879), .Y(n34437) );
  AOI32XL U36749 ( .A0(n34581), .A1(n34439), .A2(n34438), .B0(conv_2[75]), 
        .B1(n34437), .Y(n34440) );
  NAND2XL U36750 ( .A(n34440), .B(n34583), .Y(n15378) );
  OAI21XL U36751 ( .A0(n34442), .A1(n16654), .B0(n34441), .Y(n34443) );
  AOI32XL U36752 ( .A0(n34581), .A1(n34445), .A2(n34444), .B0(conv_2[450]), 
        .B1(n34443), .Y(n34446) );
  NAND2XL U36753 ( .A(n34446), .B(n34583), .Y(n15353) );
  INVXL U36754 ( .A(conv_2[90]), .Y(n34451) );
  OAI21XL U36755 ( .A0(n34448), .A1(n16655), .B0(n34447), .Y(n34449) );
  AOI32XL U36756 ( .A0(n34581), .A1(n34451), .A2(n34450), .B0(conv_2[90]), 
        .B1(n34449), .Y(n34452) );
  NAND2XL U36757 ( .A(n34452), .B(n34583), .Y(n15377) );
  AOI32XL U36758 ( .A0(n34453), .A1(n35963), .A2(n34455), .B0(n16658), .B1(
        n35963), .Y(n34454) );
  AOI32XL U36759 ( .A0(n34581), .A1(n34456), .A2(n34455), .B0(conv_2[285]), 
        .B1(n34454), .Y(n34457) );
  NAND2XL U36760 ( .A(n34457), .B(n34583), .Y(n15364) );
  OAI21XL U36761 ( .A0(n34459), .A1(n16655), .B0(n34458), .Y(n34460) );
  AOI32XL U36762 ( .A0(n34461), .A1(n34460), .A2(n34581), .B0(conv_2[225]), 
        .B1(n34460), .Y(n34462) );
  NAND2XL U36763 ( .A(n34583), .B(n34462), .Y(n15368) );
  OAI21XL U36764 ( .A0(n34463), .A1(n36042), .B0(n35986), .Y(n34464) );
  AOI32XL U36765 ( .A0(n34465), .A1(n34464), .A2(n34581), .B0(conv_2[315]), 
        .B1(n34464), .Y(n34466) );
  NAND2XL U36766 ( .A(n34583), .B(n34466), .Y(n15362) );
  NAND2XL U36767 ( .A(n34468), .B(n34467), .Y(n34470) );
  OAI21XL U36768 ( .A0(n36001), .A1(n34470), .B0(n34751), .Y(n34469) );
  AOI32XL U36769 ( .A0(n32660), .A1(n34471), .A2(n34470), .B0(conv_3[163]), 
        .B1(n34469), .Y(n34472) );
  NAND2XL U36770 ( .A(n34472), .B(n16649), .Y(n15635) );
  INVXL U36771 ( .A(conv_2[210]), .Y(n34475) );
  OAI21XL U36772 ( .A0(n34473), .A1(n16655), .B0(n35934), .Y(n34474) );
  AOI32XL U36773 ( .A0(n34476), .A1(n34475), .A2(n34581), .B0(conv_2[210]), 
        .B1(n34474), .Y(n34477) );
  NAND2XL U36774 ( .A(n34477), .B(n34583), .Y(n15369) );
  INVXL U36775 ( .A(conv_3[296]), .Y(n34483) );
  NAND2XL U36776 ( .A(n35720), .B(n34479), .Y(n34478) );
  OAI21XL U36777 ( .A0(n35720), .A1(n34479), .B0(n34478), .Y(n34481) );
  AOI211XL U36778 ( .A0(n34483), .A1(n34481), .B0(n36042), .C0(n34480), .Y(
        n34482) );
  NAND2XL U36779 ( .A(n34484), .B(n16649), .Y(n15547) );
  OAI21XL U36780 ( .A0(n34485), .A1(n16654), .B0(n36003), .Y(n34486) );
  AOI32XL U36781 ( .A0(n34581), .A1(n34486), .A2(n34525), .B0(conv_2[330]), 
        .B1(n34486), .Y(n34487) );
  NAND2XL U36782 ( .A(n34583), .B(n34487), .Y(n15361) );
  OAI21XL U36783 ( .A0(n34488), .A1(n16654), .B0(n36053), .Y(n34489) );
  AOI32XL U36784 ( .A0(n34581), .A1(n34489), .A2(n34768), .B0(conv_2[420]), 
        .B1(n34489), .Y(n34490) );
  NAND2XL U36785 ( .A(n34583), .B(n34490), .Y(n15355) );
  OAI21XL U36786 ( .A0(n34492), .A1(n16654), .B0(n34491), .Y(n34494) );
  AOI32XL U36787 ( .A0(n34581), .A1(n34494), .A2(n34493), .B0(conv_2[120]), 
        .B1(n34494), .Y(n34495) );
  NAND2XL U36788 ( .A(n34583), .B(n34495), .Y(n15375) );
  OAI21XL U36789 ( .A0(n34497), .A1(n36001), .B0(n34496), .Y(n34499) );
  AOI32XL U36790 ( .A0(n34581), .A1(n34499), .A2(n34498), .B0(conv_2[525]), 
        .B1(n34499), .Y(n34500) );
  NAND2XL U36791 ( .A(n34583), .B(n34500), .Y(n15348) );
  OAI21XL U36792 ( .A0(n34501), .A1(n16655), .B0(n36017), .Y(n34503) );
  AOI32XL U36793 ( .A0(n34581), .A1(n34503), .A2(n34502), .B0(conv_2[360]), 
        .B1(n34503), .Y(n34504) );
  NAND2XL U36794 ( .A(n34583), .B(n34504), .Y(n15359) );
  OAI21XL U36795 ( .A0(n34506), .A1(n16655), .B0(n34505), .Y(n34508) );
  AOI32XL U36796 ( .A0(n34581), .A1(n34508), .A2(n34507), .B0(conv_2[45]), 
        .B1(n34508), .Y(n34509) );
  NAND2XL U36797 ( .A(n34583), .B(n34509), .Y(n15380) );
  OAI21XL U36798 ( .A0(n34510), .A1(n16655), .B0(n35917), .Y(n34511) );
  AOI32XL U36799 ( .A0(n34581), .A1(n34511), .A2(n34706), .B0(conv_2[180]), 
        .B1(n34511), .Y(n34512) );
  NAND2XL U36800 ( .A(n34583), .B(n34512), .Y(n15371) );
  AOI22XL U36801 ( .A0(conv_3[508]), .A1(n34515), .B0(n34514), .B1(n34513), 
        .Y(n34517) );
  NAND2XL U36802 ( .A(conv_3[509]), .B(n34517), .Y(n34516) );
  OAI211XL U36803 ( .A0(conv_3[509]), .A1(n34517), .B0(n24378), .C0(n34516), 
        .Y(n34518) );
  OAI211XL U36804 ( .A0(n34520), .A1(n34519), .B0(n33468), .C0(n34518), .Y(
        n15404) );
  INVXL U36805 ( .A(conv_1[330]), .Y(n34526) );
  OAI21XL U36806 ( .A0(n34523), .A1(n16655), .B0(n35437), .Y(n34524) );
  AOI32XL U36807 ( .A0(n34769), .A1(n34526), .A2(n34525), .B0(conv_1[330]), 
        .B1(n34524), .Y(n34527) );
  NAND2XL U36808 ( .A(n34527), .B(n34773), .Y(n16133) );
  NAND2XL U36809 ( .A(n34529), .B(n34528), .Y(n34530) );
  NAND2XL U36810 ( .A(n34533), .B(n34530), .Y(n34536) );
  INVXL U36811 ( .A(n34530), .Y(n34532) );
  AOI221XL U36812 ( .A0(n34532), .A1(n36020), .B0(n34537), .B1(n16656), .C0(
        n34531), .Y(n34534) );
  AOI2BB1XL U36813 ( .A0N(n34534), .A1N(n34533), .B0(n16651), .Y(n34535) );
  OAI31XL U36814 ( .A0(n34537), .A1(n36042), .A2(n34536), .B0(n34535), .Y(
        n14947) );
  OAI21XL U36815 ( .A0(n35392), .A1(n34539), .B0(n34538), .Y(n34541) );
  AOI211XL U36816 ( .A0(n34543), .A1(n34541), .B0(n16655), .C0(n34540), .Y(
        n34542) );
  AOI2BB1XL U36817 ( .A0N(n34543), .A1N(n35395), .B0(n34542), .Y(n34545) );
  NAND2XL U36818 ( .A(n34545), .B(n34544), .Y(n16244) );
  OAI21XL U36819 ( .A0(n34548), .A1(n34547), .B0(n34546), .Y(n34550) );
  AOI211XL U36820 ( .A0(n34553), .A1(n34550), .B0(n16655), .C0(n34549), .Y(
        n34551) );
  AOI2BB1XL U36821 ( .A0N(n34553), .A1N(n34552), .B0(n34551), .Y(n34554) );
  NAND2XL U36822 ( .A(n34554), .B(n34682), .Y(n16452) );
  OAI21XL U36823 ( .A0(n34557), .A1(n34556), .B0(n34555), .Y(n34559) );
  AOI211XL U36824 ( .A0(n34561), .A1(n34559), .B0(n16655), .C0(n34558), .Y(
        n34560) );
  AOI2BB1XL U36825 ( .A0N(n34561), .A1N(n35330), .B0(n34560), .Y(n34562) );
  NAND2XL U36826 ( .A(n16652), .B(n34562), .Y(n16348) );
  NAND2XL U36827 ( .A(n34564), .B(n34563), .Y(n34566) );
  AOI211XL U36828 ( .A0(n34568), .A1(n34566), .B0(n36042), .C0(n34565), .Y(
        n34567) );
  NAND2XL U36829 ( .A(n34569), .B(n35859), .Y(n14963) );
  INVXL U36830 ( .A(conv_2[372]), .Y(n34576) );
  OAI21XL U36831 ( .A0(conv_2[371]), .A1(n34571), .B0(n34570), .Y(n34572) );
  AOI32XL U36832 ( .A0(conv_2[371]), .A1(n34572), .A2(n34571), .B0(n34570), 
        .B1(n34572), .Y(n34574) );
  AOI211XL U36833 ( .A0(n34576), .A1(n34574), .B0(n36001), .C0(n34573), .Y(
        n34575) );
  NAND2XL U36834 ( .A(n34577), .B(n35859), .Y(n14956) );
  OAI21XL U36835 ( .A0(n34578), .A1(n16655), .B0(n34631), .Y(n34580) );
  AOI32XL U36836 ( .A0(n34581), .A1(n34580), .A2(n34579), .B0(conv_2[150]), 
        .B1(n34580), .Y(n34582) );
  NAND2XL U36837 ( .A(n34583), .B(n34582), .Y(n15373) );
  INVXL U36838 ( .A(conv_2[177]), .Y(n34590) );
  NAND2XL U36839 ( .A(n29831), .B(n34585), .Y(n34584) );
  OAI21XL U36840 ( .A0(n29831), .A1(n34585), .B0(n34584), .Y(n34587) );
  AOI211XL U36841 ( .A0(n34590), .A1(n34587), .B0(n16655), .C0(n34586), .Y(
        n34588) );
  NAND2XL U36842 ( .A(n34591), .B(n34735), .Y(n15086) );
  OAI211XL U36843 ( .A0(conv_2[179]), .A1(n34596), .B0(n16657), .C0(n34595), 
        .Y(n34597) );
  OAI21XL U36844 ( .A0(n34603), .A1(n34389), .B0(n34601), .Y(n34602) );
  AOI32XL U36845 ( .A0(n33788), .A1(n34604), .A2(n34603), .B0(conv_2[261]), 
        .B1(n34602), .Y(n34605) );
  NAND2XL U36846 ( .A(n34605), .B(n34735), .Y(n15032) );
  NAND2BXL U36847 ( .AN(n34607), .B(n34606), .Y(n34609) );
  AOI211XL U36848 ( .A0(n34611), .A1(n34609), .B0(n16655), .C0(n34608), .Y(
        n34610) );
  NAND2XL U36849 ( .A(n34612), .B(n35566), .Y(n15846) );
  NAND2XL U36850 ( .A(n34614), .B(n34613), .Y(n34616) );
  NAND2XL U36851 ( .A(n34616), .B(n34615), .Y(n34618) );
  AOI211XL U36852 ( .A0(n34620), .A1(n34618), .B0(n16655), .C0(n34617), .Y(
        n34619) );
  NAND2XL U36853 ( .A(n34622), .B(n34621), .Y(n15302) );
  INVXL U36854 ( .A(conv_2[160]), .Y(n34632) );
  AOI32XL U36855 ( .A0(n34627), .A1(n34626), .A2(n34625), .B0(n34624), .B1(
        n34623), .Y(n34629) );
  AOI211XL U36856 ( .A0(n34632), .A1(n34629), .B0(n16655), .C0(n34628), .Y(
        n34630) );
  NAND2XL U36857 ( .A(n34633), .B(n35859), .Y(n15098) );
  AOI32XL U36858 ( .A0(conv_2[398]), .A1(n34636), .A2(n34635), .B0(n34634), 
        .B1(n34636), .Y(n34638) );
  AOI211XL U36859 ( .A0(n34640), .A1(n34638), .B0(n16655), .C0(n34637), .Y(
        n34639) );
  AOI2BB1XL U36860 ( .A0N(n34640), .A1N(n36031), .B0(n34639), .Y(n34641) );
  NAND2XL U36861 ( .A(n34641), .B(n35859), .Y(n14939) );
  NAND2XL U36862 ( .A(n34643), .B(n34642), .Y(n34645) );
  AOI211XL U36863 ( .A0(n34647), .A1(n34645), .B0(n16655), .C0(n34644), .Y(
        n34646) );
  AOI2BB1XL U36864 ( .A0N(n34647), .A1N(n35894), .B0(n34646), .Y(n34648) );
  NAND2XL U36865 ( .A(n34648), .B(n35859), .Y(n15127) );
  AOI32XL U36866 ( .A0(conv_3[221]), .A1(n34649), .A2(n35667), .B0(n35660), 
        .B1(n35668), .Y(n34651) );
  AOI211XL U36867 ( .A0(n34653), .A1(n34651), .B0(n16655), .C0(n34650), .Y(
        n34652) );
  AOI2BB1XL U36868 ( .A0N(n34653), .A1N(n35665), .B0(n34652), .Y(n34654) );
  NAND2XL U36869 ( .A(n34654), .B(n35588), .Y(n15596) );
  INVXL U36870 ( .A(conv_3[203]), .Y(n34660) );
  NAND2XL U36871 ( .A(n35653), .B(n34656), .Y(n34655) );
  OAI21XL U36872 ( .A0(n35653), .A1(n34656), .B0(n34655), .Y(n34658) );
  AOI211XL U36873 ( .A0(n34660), .A1(n34658), .B0(n16655), .C0(n34657), .Y(
        n34659) );
  AOI2BB1XL U36874 ( .A0N(n34660), .A1N(n35646), .B0(n34659), .Y(n34661) );
  NAND2XL U36875 ( .A(n34661), .B(n35588), .Y(n15610) );
  AOI22XL U36876 ( .A0(conv_2[493]), .A1(n34664), .B0(n34663), .B1(n34662), 
        .Y(n34667) );
  NAND2XL U36877 ( .A(conv_2[494]), .B(n34667), .Y(n34665) );
  OAI211XL U36878 ( .A0(conv_2[494]), .A1(n34667), .B0(n34666), .C0(n34665), 
        .Y(n34668) );
  OAI211XL U36879 ( .A0(n34789), .A1(n34670), .B0(n34669), .C0(n34668), .Y(
        n14874) );
  NAND2XL U36880 ( .A(n34776), .B(n34775), .Y(n34774) );
  INVXL U36881 ( .A(conv_1[418]), .Y(n34778) );
  OAI32XL U36882 ( .A0(conv_1[418]), .A1(n34776), .A2(n34775), .B0(n34774), 
        .B1(n34778), .Y(n34673) );
  NAND2XL U36883 ( .A(conv_1[419]), .B(n34673), .Y(n34672) );
  OAI211XL U36884 ( .A0(conv_1[419]), .A1(n34673), .B0(n32181), .C0(n34672), 
        .Y(n34674) );
  OAI211XL U36885 ( .A0(n34676), .A1(n34675), .B0(n34696), .C0(n34674), .Y(
        n16044) );
  NAND2XL U36886 ( .A(n34678), .B(n34677), .Y(n34680) );
  OAI21XL U36887 ( .A0(n16655), .A1(n34680), .B0(n35395), .Y(n34679) );
  AOI32XL U36888 ( .A0(n36020), .A1(n34681), .A2(n34680), .B0(conv_1[223]), 
        .B1(n34679), .Y(n34683) );
  NAND2XL U36889 ( .A(n34683), .B(n34682), .Y(n16240) );
  NAND2XL U36890 ( .A(n34685), .B(n34684), .Y(n34687) );
  OAI21XL U36891 ( .A0(n16655), .A1(n34687), .B0(n35346), .Y(n34686) );
  AOI32XL U36892 ( .A0(n33778), .A1(n34688), .A2(n34687), .B0(conv_1[178]), 
        .B1(n34686), .Y(n34690) );
  NAND2XL U36893 ( .A(n34690), .B(n34689), .Y(n16285) );
  NAND2XL U36894 ( .A(n34692), .B(n34691), .Y(n34694) );
  OAI21XL U36895 ( .A0(n16655), .A1(n34694), .B0(n35477), .Y(n34693) );
  AOI32XL U36896 ( .A0(n30090), .A1(n34695), .A2(n34694), .B0(conv_1[403]), 
        .B1(n34693), .Y(n34697) );
  NAND2XL U36897 ( .A(n34697), .B(n34696), .Y(n16060) );
  OAI21XL U36898 ( .A0(n34698), .A1(n16655), .B0(n35598), .Y(n34700) );
  AOI32XL U36899 ( .A0(n34742), .A1(n34700), .A2(n34699), .B0(conv_3[60]), 
        .B1(n34700), .Y(n34701) );
  NAND2XL U36900 ( .A(n34755), .B(n34701), .Y(n15919) );
  OAI21XL U36901 ( .A0(n34705), .A1(n16655), .B0(n34704), .Y(n34707) );
  AOI32XL U36902 ( .A0(n34742), .A1(n34707), .A2(n34706), .B0(conv_3[180]), 
        .B1(n34707), .Y(n34708) );
  NAND2XL U36903 ( .A(n34755), .B(n34708), .Y(n15911) );
  OAI21XL U36904 ( .A0(n34710), .A1(n16655), .B0(n34709), .Y(n34712) );
  AOI32XL U36905 ( .A0(n34742), .A1(n34712), .A2(n34711), .B0(conv_3[270]), 
        .B1(n34712), .Y(n34713) );
  NAND2XL U36906 ( .A(n34755), .B(n34713), .Y(n15905) );
  OAI21XL U36907 ( .A0(n34716), .A1(n16654), .B0(n35330), .Y(n34718) );
  AOI32XL U36908 ( .A0(n34769), .A1(n34718), .A2(n34717), .B0(conv_1[105]), 
        .B1(n34718), .Y(n34719) );
  NAND2XL U36909 ( .A(n34773), .B(n34719), .Y(n16358) );
  OAI21XL U36910 ( .A0(n34720), .A1(n16654), .B0(n35576), .Y(n34722) );
  AOI32XL U36911 ( .A0(n34742), .A1(n34722), .A2(n34721), .B0(conv_3[15]), 
        .B1(n34722), .Y(n34723) );
  NAND2XL U36912 ( .A(n34755), .B(n34723), .Y(n15922) );
  NAND2XL U36913 ( .A(n34725), .B(n34724), .Y(n34727) );
  OAI21XL U36914 ( .A0(n16655), .A1(n34727), .B0(n35846), .Y(n34726) );
  AOI32XL U36915 ( .A0(n33778), .A1(n34728), .A2(n34727), .B0(conv_2[73]), 
        .B1(n34726), .Y(n34729) );
  NAND2XL U36916 ( .A(n34729), .B(n34735), .Y(n15155) );
  NAND2XL U36917 ( .A(n34731), .B(n34730), .Y(n34733) );
  OAI21XL U36918 ( .A0(n16655), .A1(n34733), .B0(n36070), .Y(n34732) );
  NAND2XL U36919 ( .A(n34736), .B(n34735), .Y(n14905) );
  INVXL U36920 ( .A(conv_3[135]), .Y(n34741) );
  AOI32XL U36921 ( .A0(n34738), .A1(n34737), .A2(n34740), .B0(n16655), .B1(
        n34737), .Y(n34739) );
  AOI32XL U36922 ( .A0(n34742), .A1(n34741), .A2(n34740), .B0(conv_3[135]), 
        .B1(n34739), .Y(n34743) );
  NAND2XL U36923 ( .A(n34743), .B(n34755), .Y(n15914) );
  NAND2XL U36924 ( .A(n34745), .B(n34744), .Y(n34748) );
  OAI21XL U36925 ( .A0(n16655), .A1(n34748), .B0(n34746), .Y(n34747) );
  AOI32XL U36926 ( .A0(n32656), .A1(n34749), .A2(n34748), .B0(conv_3[358]), 
        .B1(n34747), .Y(n34750) );
  NAND2XL U36927 ( .A(n34750), .B(n35588), .Y(n15505) );
  INVXL U36928 ( .A(conv_3[150]), .Y(n34754) );
  OAI21XL U36929 ( .A0(n16655), .A1(n34753), .B0(n34751), .Y(n34752) );
  NAND2XL U36930 ( .A(n34756), .B(n34755), .Y(n15913) );
  INVXL U36931 ( .A(conv_3[133]), .Y(n34781) );
  OAI21XL U36932 ( .A0(n34784), .A1(n34783), .B0(n34782), .Y(n34759) );
  NAND2XL U36933 ( .A(conv_3[133]), .B(n34759), .Y(n34758) );
  OAI211XL U36934 ( .A0(conv_3[133]), .A1(n34759), .B0(n34028), .C0(n34758), 
        .Y(n34760) );
  OAI211XL U36935 ( .A0(n35626), .A1(n34781), .B0(n16649), .C0(n34760), .Y(
        n15655) );
  INVXL U36936 ( .A(conv_1[345]), .Y(n34761) );
  OAI2BB1XL U36937 ( .A0N(n34769), .A1N(n34762), .B0(n34761), .Y(n34765) );
  AOI32XL U36938 ( .A0(n16656), .A1(n34765), .A2(n34764), .B0(n34763), .B1(
        n34765), .Y(n34766) );
  NAND2XL U36939 ( .A(n34773), .B(n34766), .Y(n16118) );
  INVXL U36940 ( .A(conv_1[420]), .Y(n34767) );
  OAI2BB1XL U36941 ( .A0N(n34769), .A1N(n34768), .B0(n34767), .Y(n34771) );
  AOI32XL U36942 ( .A0(n33822), .A1(n34771), .A2(n34770), .B0(n35510), .B1(
        n34771), .Y(n34772) );
  NAND2XL U36943 ( .A(n34773), .B(n34772), .Y(n16043) );
  OAI2BB2XL U36944 ( .B0(conv_1[418]), .B1(n34777), .A0N(conv_1[418]), .A1N(
        n34777), .Y(n34779) );
  OAI22XL U36945 ( .A0(n36001), .A1(n34779), .B0(n35487), .B1(n34778), .Y(
        n34780) );
  OR2XL U36946 ( .A(n35549), .B(n34780), .Y(n16045) );
  OAI211XL U36947 ( .A0(conv_3[134]), .A1(n34786), .B0(n32611), .C0(n34785), 
        .Y(n34787) );
  OAI211XL U36948 ( .A0(n34789), .A1(n34788), .B0(n16649), .C0(n34787), .Y(
        n15654) );
  AOI2BB2XL U36950 ( .B0(n34798), .B1(n34797), .A0N(pool[6]), .A1N(n34798), 
        .Y(N29222) );
  AOI2BB2XL U36951 ( .B0(n34806), .B1(n34805), .A0N(n34804), .A1N(n34806), .Y(
        N29228) );
  AOI2BB2XL U36952 ( .B0(n34808), .B1(n34807), .A0N(pool[16]), .A1N(n34808), 
        .Y(N29232) );
  AOI2BB2XL U36953 ( .B0(n34821), .B1(n34820), .A0N(n34819), .A1N(n34821), .Y(
        N29243) );
  OAI22XL U36954 ( .A0(n34823), .A1(n28349), .B0(n34822), .B1(n26621), .Y(
        n34833) );
  AOI22XL U36955 ( .A0(n16670), .A1(n34825), .B0(n16664), .B1(n34824), .Y(
        n34830) );
  AOI22XL U36956 ( .A0(n35130), .A1(n34828), .B0(n34827), .B1(n34826), .Y(
        n34829) );
  OAI211XL U36957 ( .A0(n35135), .A1(n34831), .B0(n34830), .C0(n34829), .Y(
        n34832) );
  OAI2BB2XL U36958 ( .B0(n34839), .B1(n34834), .A0N(pool[30]), .A1N(n34839), 
        .Y(N29246) );
  AOI22XL U36959 ( .A0(n35195), .A1(n34846), .B0(n35234), .B1(n34845), .Y(
        n34850) );
  AOI22XL U36960 ( .A0(n35236), .A1(n34848), .B0(n34847), .B1(n35231), .Y(
        n34849) );
  OAI211XL U36961 ( .A0(n34851), .A1(n35198), .B0(n34850), .C0(n34849), .Y(
        n34855) );
  OAI22XL U36962 ( .A0(N18471), .A1(n34853), .B0(n34852), .B1(n35135), .Y(
        n34854) );
  OAI2BB2XL U36963 ( .B0(n34860), .B1(n34856), .A0N(pool[40]), .A1N(n34860), 
        .Y(N29256) );
  AOI2BB2XL U36964 ( .B0(n34864), .B1(n34863), .A0N(pool[46]), .A1N(n34864), 
        .Y(N29262) );
  AOI2BB2XL U36965 ( .B0(n34881), .B1(n34885), .A0N(n34885), .A1N(pool[61]), 
        .Y(N29277) );
  AOI2BB2XL U36966 ( .B0(n34884), .B1(n34883), .A0N(n34882), .A1N(n34884), .Y(
        N29278) );
  AOI2BB2XL U36967 ( .B0(n34886), .B1(n34885), .A0N(n34885), .A1N(pool[63]), 
        .Y(N29279) );
  AOI2BB2XL U36968 ( .B0(n34896), .B1(n34895), .A0N(n34894), .A1N(n34896), .Y(
        N29288) );
  AOI2BB2XL U36969 ( .B0(n34901), .B1(n34900), .A0N(n34899), .A1N(n34901), .Y(
        N29293) );
  AOI22XL U36970 ( .A0(n28528), .A1(n34904), .B0(n34903), .B1(n34902), .Y(
        n34909) );
  AOI22XL U36971 ( .A0(n35236), .A1(n34907), .B0(n34906), .B1(n34905), .Y(
        n34908) );
  OAI211XL U36972 ( .A0(n34910), .A1(n16672), .B0(n34909), .C0(n34908), .Y(
        n34919) );
  AOI22XL U36973 ( .A0(n19179), .A1(n34912), .B0(n16671), .B1(n34911), .Y(
        n34916) );
  AOI22XL U36974 ( .A0(n35195), .A1(n34914), .B0(n18197), .B1(n34913), .Y(
        n34915) );
  OAI211XL U36975 ( .A0(n34917), .A1(n35159), .B0(n34916), .C0(n34915), .Y(
        n34918) );
  AOI211XL U36976 ( .A0(n34921), .A1(n34920), .B0(n34919), .C0(n34918), .Y(
        n34923) );
  AOI2BB2XL U36977 ( .B0(n34926), .B1(n34925), .A0N(n34924), .A1N(n34926), .Y(
        N29298) );
  OAI2BB2XL U36978 ( .B0(N18471), .B1(n34928), .A0N(n34927), .A1N(n16700), .Y(
        n34937) );
  AOI22XL U36979 ( .A0(n35195), .A1(n34930), .B0(n35236), .B1(n34929), .Y(
        n34934) );
  AOI22XL U36980 ( .A0(n35234), .A1(n34932), .B0(n34931), .B1(n35231), .Y(
        n34933) );
  OAI211XL U36981 ( .A0(n34935), .A1(n35198), .B0(n34934), .C0(n34933), .Y(
        n34936) );
  OAI2BB2XL U36982 ( .B0(n34940), .B1(n34938), .A0N(pool[85]), .A1N(n34940), 
        .Y(N29301) );
  AOI22XL U36983 ( .A0(n34952), .A1(n34951), .B0(n34950), .B1(n34949), .Y(
        n34957) );
  AOI22XL U36984 ( .A0(n16667), .A1(n34955), .B0(n34954), .B1(n34953), .Y(
        n34956) );
  OAI211XL U36985 ( .A0(n34959), .A1(n34958), .B0(n34957), .C0(n34956), .Y(
        n34971) );
  AOI22XL U36986 ( .A0(n28528), .A1(n34965), .B0(n35234), .B1(n34964), .Y(
        n34966) );
  OAI211XL U36987 ( .A0(n34969), .A1(n34968), .B0(n34967), .C0(n34966), .Y(
        n34970) );
  AOI211XL U36988 ( .A0(n28465), .A1(n34972), .B0(n34971), .C0(n34970), .Y(
        n34974) );
  INVXL U36989 ( .A(pool[95]), .Y(n34973) );
  OAI22XL U36990 ( .A0(n34983), .A1(n34982), .B0(n35240), .B1(n34981), .Y(
        n34991) );
  AOI22XL U36991 ( .A0(n16667), .A1(n35232), .B0(n34984), .B1(n35233), .Y(
        n34988) );
  AOI22XL U36992 ( .A0(n16665), .A1(n34986), .B0(n16671), .B1(n34985), .Y(
        n34987) );
  OAI211XL U36993 ( .A0(n34989), .A1(n35242), .B0(n34988), .C0(n34987), .Y(
        n34990) );
  AOI211XL U36994 ( .A0(n34992), .A1(n35235), .B0(n34991), .C0(n34990), .Y(
        n34994) );
  NAND2XL U36995 ( .A(n35010), .B(pool[105]), .Y(n35002) );
  OAI2BB1XL U36996 ( .A0N(n35003), .A1N(n35006), .B0(n35002), .Y(N29321) );
  AOI2BB2XL U36997 ( .B0(n35022), .B1(n35021), .A0N(n35020), .A1N(n35022), .Y(
        N29338) );
  OAI22XL U36998 ( .A0(n35030), .A1(n35196), .B0(n35029), .B1(n18208), .Y(
        n35039) );
  AOI22XL U36999 ( .A0(n35181), .A1(n35032), .B0(n16664), .B1(n35031), .Y(
        n35036) );
  AOI2BB2XL U37000 ( .B0(n35207), .B1(n35034), .A0N(n35198), .A1N(n35033), .Y(
        n35035) );
  OAI211XL U37001 ( .A0(n35135), .A1(n35037), .B0(n35036), .C0(n35035), .Y(
        n35038) );
  AOI211XL U37002 ( .A0(n35195), .A1(n35040), .B0(n35039), .C0(n35038), .Y(
        n35215) );
  OAI22XL U37003 ( .A0(n35042), .A1(n35202), .B0(n35041), .B1(n18208), .Y(
        n35051) );
  AOI22XL U37004 ( .A0(n35234), .A1(n35044), .B0(n16664), .B1(n35043), .Y(
        n35048) );
  AOI22XL U37005 ( .A0(n16660), .A1(n35046), .B0(n35207), .B1(n35045), .Y(
        n35047) );
  OAI211XL U37006 ( .A0(n35135), .A1(n35049), .B0(n35048), .C0(n35047), .Y(
        n35050) );
  AOI211XL U37007 ( .A0(n35195), .A1(n35052), .B0(n35051), .C0(n35050), .Y(
        n35216) );
  NAND2XL U37008 ( .A(n35215), .B(n35216), .Y(n35125) );
  AOI2BB2XL U37009 ( .B0(n35207), .B1(n35054), .A0N(n35196), .A1N(n35053), .Y(
        n35063) );
  OAI22XL U37010 ( .A0(n35056), .A1(n35200), .B0(n35055), .B1(n35202), .Y(
        n35060) );
  OAI22XL U37011 ( .A0(n35058), .A1(n18208), .B0(n35057), .B1(n35198), .Y(
        n35059) );
  AOI211XL U37012 ( .A0(n35195), .A1(n35061), .B0(n35060), .C0(n35059), .Y(
        n35062) );
  OAI211XL U37013 ( .A0(n35135), .A1(n35064), .B0(n35063), .C0(n35062), .Y(
        n35213) );
  AOI2BB2XL U37014 ( .B0(n16664), .B1(n35066), .A0N(n35196), .A1N(n35065), .Y(
        n35075) );
  OAI22XL U37015 ( .A0(n35068), .A1(n35202), .B0(n35067), .B1(n18208), .Y(
        n35072) );
  OAI2BB2XL U37016 ( .B0(n35184), .B1(n35070), .A0N(n35069), .A1N(n16660), .Y(
        n35071) );
  AOI211XL U37017 ( .A0(n35195), .A1(n35073), .B0(n35072), .C0(n35071), .Y(
        n35074) );
  OAI211XL U37018 ( .A0(n35241), .A1(n35076), .B0(n35075), .C0(n35074), .Y(
        n35211) );
  OAI22XL U37019 ( .A0(n35078), .A1(n35200), .B0(n35077), .B1(n35196), .Y(
        n35087) );
  AOI22XL U37020 ( .A0(n35181), .A1(n35080), .B0(n35236), .B1(n35079), .Y(
        n35084) );
  AOI2BB2XL U37021 ( .B0(n35195), .B1(n35082), .A0N(n35184), .A1N(n35081), .Y(
        n35083) );
  OAI211XL U37022 ( .A0(n35085), .A1(n35198), .B0(n35084), .C0(n35083), .Y(
        n35086) );
  AOI211XL U37023 ( .A0(n28465), .A1(n35088), .B0(n35087), .C0(n35086), .Y(
        n35212) );
  OAI22XL U37024 ( .A0(n35184), .A1(n35090), .B0(n35089), .B1(n35200), .Y(
        n35099) );
  AOI22XL U37025 ( .A0(n35195), .A1(n35092), .B0(n35236), .B1(n35091), .Y(
        n35096) );
  AOI22XL U37026 ( .A0(n35181), .A1(n35094), .B0(n35234), .B1(n35093), .Y(
        n35095) );
  OAI211XL U37027 ( .A0(n35135), .A1(n35097), .B0(n35096), .C0(n35095), .Y(
        n35098) );
  AOI211XL U37028 ( .A0(n16660), .A1(n35100), .B0(n35099), .C0(n35098), .Y(
        n35220) );
  AOI22XL U37029 ( .A0(n35236), .A1(n35102), .B0(n16660), .B1(n35101), .Y(
        n35106) );
  AOI2BB2XL U37030 ( .B0(n35231), .B1(n35104), .A0N(n35196), .A1N(n35103), .Y(
        n35105) );
  OAI211XL U37031 ( .A0(n35107), .A1(n35239), .B0(n35106), .C0(n35105), .Y(
        n35111) );
  OAI22XL U37032 ( .A0(n35109), .A1(n35159), .B0(n35135), .B1(n35108), .Y(
        n35110) );
  OAI22XL U37033 ( .A0(n35113), .A1(n35198), .B0(n35112), .B1(n35200), .Y(
        n35122) );
  AOI22XL U37034 ( .A0(n35195), .A1(n35115), .B0(n35207), .B1(n35114), .Y(
        n35119) );
  AOI22XL U37035 ( .A0(n35236), .A1(n35117), .B0(n35234), .B1(n35116), .Y(
        n35118) );
  OAI211XL U37036 ( .A0(n35135), .A1(n35120), .B0(n35119), .C0(n35118), .Y(
        n35121) );
  AOI211XL U37037 ( .A0(n35181), .A1(n35123), .B0(n35122), .C0(n35121), .Y(
        n35219) );
  NAND4XL U37038 ( .A(n35212), .B(n35220), .C(n35253), .D(n35219), .Y(n35124)
         );
  AOI2BB2XL U37039 ( .B0(n35236), .B1(n35127), .A0N(n35239), .A1N(n35126), .Y(
        n35132) );
  AOI22XL U37040 ( .A0(n35130), .A1(n35129), .B0(n16660), .B1(n35128), .Y(
        n35131) );
  OAI211XL U37041 ( .A0(n35143), .A1(n35133), .B0(n35132), .C0(n35131), .Y(
        n35138) );
  OAI22XL U37042 ( .A0(n35136), .A1(n35159), .B0(n35135), .B1(n35134), .Y(
        n35137) );
  INVXL U37043 ( .A(pool[132]), .Y(n35249) );
  AOI22XL U37044 ( .A0(n35236), .A1(n35140), .B0(n35234), .B1(n35139), .Y(
        n35150) );
  OAI22XL U37045 ( .A0(n35143), .A1(n35142), .B0(n35141), .B1(n35198), .Y(
        n35147) );
  OAI22XL U37046 ( .A0(N18471), .A1(n35145), .B0(n35144), .B1(n35135), .Y(
        n35146) );
  AOI211XL U37047 ( .A0(n35195), .A1(n35148), .B0(n35147), .C0(n35146), .Y(
        n35149) );
  NAND2XL U37048 ( .A(n35150), .B(n35149), .Y(n35248) );
  AOI22XL U37049 ( .A0(n35195), .A1(n35152), .B0(n16660), .B1(n35151), .Y(
        n35156) );
  AOI22XL U37050 ( .A0(n35236), .A1(n35154), .B0(n35231), .B1(n35153), .Y(
        n35155) );
  OAI211XL U37051 ( .A0(n35157), .A1(n35196), .B0(n35156), .C0(n35155), .Y(
        n35162) );
  OAI22XL U37052 ( .A0(n35160), .A1(n35159), .B0(n35135), .B1(n35158), .Y(
        n35161) );
  AOI222XL U37053 ( .A0(pool[130]), .A1(pool[131]), .B0(pool[130]), .B1(n35247), .C0(pool[131]), .C1(n35247), .Y(n35163) );
  AOI222XL U37054 ( .A0(n35249), .A1(n35248), .B0(n35249), .B1(n35163), .C0(
        n35248), .C1(n35163), .Y(n35164) );
  AOI222XL U37055 ( .A0(n35251), .A1(pool[133]), .B0(n35251), .B1(n35164), 
        .C0(pool[133]), .C1(n35164), .Y(n35165) );
  AOI22XL U37056 ( .A0(n35195), .A1(n35168), .B0(n16660), .B1(n35167), .Y(
        n35177) );
  OAI2BB2XL U37057 ( .B0(n35170), .B1(n35196), .A0N(n35207), .A1N(n35169), .Y(
        n35174) );
  OAI22XL U37058 ( .A0(n35172), .A1(n18208), .B0(n35171), .B1(n35200), .Y(
        n35173) );
  AOI211XL U37059 ( .A0(n28465), .A1(n35175), .B0(n35174), .C0(n35173), .Y(
        n35176) );
  OAI211XL U37060 ( .A0(n35178), .A1(n35202), .B0(n35177), .C0(n35176), .Y(
        n35225) );
  AOI22XL U37061 ( .A0(n35181), .A1(n35180), .B0(n35195), .B1(n35179), .Y(
        n35191) );
  OAI22XL U37062 ( .A0(n35184), .A1(n35183), .B0(n35182), .B1(n35200), .Y(
        n35188) );
  OAI2BB2XL U37063 ( .B0(n35186), .B1(n35196), .A0N(n35185), .A1N(n16660), .Y(
        n35187) );
  AOI211XL U37064 ( .A0(n35236), .A1(n35189), .B0(n35188), .C0(n35187), .Y(
        n35190) );
  OAI211XL U37065 ( .A0(n35135), .A1(n35192), .B0(n35191), .C0(n35190), .Y(
        n35221) );
  AOI22XL U37066 ( .A0(n35195), .A1(n35194), .B0(n35236), .B1(n35193), .Y(
        n35209) );
  OAI22XL U37067 ( .A0(n35199), .A1(n35198), .B0(n35197), .B1(n35196), .Y(
        n35205) );
  OAI22XL U37068 ( .A0(n35203), .A1(n35202), .B0(n35201), .B1(n35200), .Y(
        n35204) );
  AOI211XL U37069 ( .A0(n35207), .A1(n35206), .B0(n35205), .C0(n35204), .Y(
        n35208) );
  OAI211XL U37070 ( .A0(n35135), .A1(n35210), .B0(n35209), .C0(n35208), .Y(
        n35214) );
  NOR3XL U37071 ( .A(pool[134]), .B(n35221), .C(n35214), .Y(n35224) );
  NAND2BXL U37072 ( .AN(n35212), .B(n35211), .Y(n35218) );
  NAND4BBXL U37073 ( .AN(n35216), .BN(n35215), .C(n35214), .D(n35213), .Y(
        n35217) );
  NOR4XL U37074 ( .A(n35220), .B(n35219), .C(n35218), .D(n35217), .Y(n35222)
         );
  NAND4BXL U37075 ( .AN(n35253), .B(pool[134]), .C(n35222), .D(n35221), .Y(
        n35223) );
  AOI22XL U37076 ( .A0(n16660), .A1(n35232), .B0(n35231), .B1(n35230), .Y(
        n35238) );
  AOI22XL U37077 ( .A0(n35236), .A1(n35235), .B0(n35234), .B1(n35233), .Y(
        n35237) );
  OAI211XL U37078 ( .A0(n35240), .A1(n35239), .B0(n35238), .C0(n35237), .Y(
        n35245) );
  OAI22XL U37079 ( .A0(N18471), .A1(n35243), .B0(n35242), .B1(n35241), .Y(
        n35244) );
  OAI2BB2XL U37080 ( .B0(n35250), .B1(n35246), .A0N(pool[130]), .A1N(n35250), 
        .Y(N29346) );
  OAI21XL U37081 ( .A0(n36244), .A1(n35255), .B0(n35265), .Y(n35257) );
  OAI2BB2XL U37082 ( .B0(n35258), .B1(n35257), .A0N(n35256), .A1N(N29500), .Y(
        n16643) );
  AOI31XL U37083 ( .A0(n35265), .A1(n16669), .A2(n35262), .B0(n35264), .Y(
        n35263) );
  OAI2BB1XL U37084 ( .A0N(N29497), .A1N(n35267), .B0(n35263), .Y(n16640) );
  AOI31XL U37085 ( .A0(n35265), .A1(n19902), .A2(n22612), .B0(n35264), .Y(
        n35266) );
  OAI2BB1XL U37086 ( .A0N(N29496), .A1N(n35267), .B0(n35266), .Y(n16639) );
  OAI2BB2XL U37087 ( .B0(n35272), .B1(n35271), .A0N(n35270), .A1N(conv_1[1]), 
        .Y(intadd_2_CI) );
  AOI2BB1XL U37088 ( .A0N(n35275), .A1N(n35274), .B0(n35273), .Y(n35276) );
  OAI2BB2XL U37089 ( .B0(conv_1[25]), .B1(n35276), .A0N(conv_1[25]), .A1N(
        n35276), .Y(n35279) );
  OAI22XL U37090 ( .A0(n36009), .A1(n35279), .B0(n35278), .B1(n35277), .Y(
        n35280) );
  OR2XL U37091 ( .A(n35549), .B(n35280), .Y(n16438) );
  AOI2BB1XL U37092 ( .A0N(n35296), .A1N(n35282), .B0(n35281), .Y(n35283) );
  OAI2BB2XL U37093 ( .B0(conv_1[36]), .B1(n35283), .A0N(conv_1[36]), .A1N(
        n35283), .Y(n35285) );
  OAI22XL U37094 ( .A0(n16654), .A1(n35285), .B0(n35302), .B1(n35284), .Y(
        n35286) );
  OR2XL U37095 ( .A(n35549), .B(n35286), .Y(n16427) );
  AOI21XL U37096 ( .A0(n35289), .A1(n35288), .B0(n35287), .Y(n35290) );
  OAI2BB2XL U37097 ( .B0(conv_1[37]), .B1(n35290), .A0N(conv_1[37]), .A1N(
        n35290), .Y(n35292) );
  OAI22XL U37098 ( .A0(n16658), .A1(n35292), .B0(n35302), .B1(n35291), .Y(
        n35293) );
  OR2XL U37099 ( .A(n35549), .B(n35293), .Y(n16426) );
  AOI2BB1XL U37100 ( .A0N(n35296), .A1N(n35295), .B0(n35294), .Y(n35297) );
  OAI2BB2XL U37101 ( .B0(conv_1[40]), .B1(n35297), .A0N(conv_1[40]), .A1N(
        n35297), .Y(n35299) );
  OAI22XL U37102 ( .A0(n36009), .A1(n35299), .B0(n35302), .B1(n35298), .Y(
        n35300) );
  OR2XL U37103 ( .A(n35549), .B(n35300), .Y(n16423) );
  AOI32XL U37104 ( .A0(n35303), .A1(n35302), .A2(n35301), .B0(n36009), .B1(
        n35302), .Y(n35306) );
  AOI21XL U37105 ( .A0(n35309), .A1(n35308), .B0(n35307), .Y(n35310) );
  OAI2BB2XL U37106 ( .B0(conv_1[54]), .B1(n35310), .A0N(conv_1[54]), .A1N(
        n35310), .Y(n35312) );
  OAI22XL U37107 ( .A0(n34389), .A1(n35312), .B0(n35319), .B1(n35311), .Y(
        n35313) );
  AOI2BB1XL U37108 ( .A0N(n35316), .A1N(n35315), .B0(n35314), .Y(n35317) );
  OAI2BB2XL U37109 ( .B0(conv_1[55]), .B1(n35317), .A0N(conv_1[55]), .A1N(
        n35317), .Y(n35320) );
  OAI22XL U37110 ( .A0(n36042), .A1(n35320), .B0(n35319), .B1(n35318), .Y(
        n35321) );
  OR2XL U37111 ( .A(n35549), .B(n35321), .Y(n16408) );
  AOI21XL U37112 ( .A0(n35324), .A1(n35323), .B0(n35322), .Y(n35325) );
  OAI2BB2XL U37113 ( .B0(conv_1[67]), .B1(n35325), .A0N(conv_1[67]), .A1N(
        n35325), .Y(n35328) );
  OAI22XL U37114 ( .A0(n16654), .A1(n35328), .B0(n35327), .B1(n35326), .Y(
        n35329) );
  OR2XL U37115 ( .A(n35549), .B(n35329), .Y(n16396) );
  AOI32XL U37116 ( .A0(n35331), .A1(n35330), .A2(n35332), .B0(n36042), .B1(
        n35330), .Y(n35335) );
  AOI31XL U37117 ( .A0(n36020), .A1(n35333), .A2(n35332), .B0(n35549), .Y(
        n35334) );
  OAI2BB1XL U37118 ( .A0N(conv_1[116]), .A1N(n35335), .B0(n35334), .Y(n16347)
         );
  AOI2BB1XL U37119 ( .A0N(n35339), .A1N(n35338), .B0(n35337), .Y(n35340) );
  OAI2BB2XL U37120 ( .B0(conv_1[142]), .B1(n35340), .A0N(conv_1[142]), .A1N(
        n35340), .Y(n35342) );
  OAI2BB2XL U37121 ( .B0(n16654), .B1(n35342), .A0N(n35341), .A1N(conv_1[142]), 
        .Y(n35343) );
  OR2XL U37122 ( .A(n35549), .B(n35343), .Y(n16321) );
  INVXL U37123 ( .A(n35344), .Y(n35345) );
  AOI32XL U37124 ( .A0(n35347), .A1(n35346), .A2(n35345), .B0(n36001), .B1(
        n35346), .Y(n35350) );
  AOI31XL U37125 ( .A0(n36020), .A1(n35348), .A2(n35347), .B0(n35549), .Y(
        n35349) );
  OAI2BB1XL U37126 ( .A0N(conv_1[170]), .A1N(n35350), .B0(n35349), .Y(n16293)
         );
  AOI2BB1XL U37127 ( .A0N(n35365), .A1N(n35352), .B0(n35351), .Y(n35353) );
  OAI2BB2XL U37128 ( .B0(conv_1[186]), .B1(n35353), .A0N(conv_1[186]), .A1N(
        n35353), .Y(n35355) );
  OAI22XL U37129 ( .A0(n36009), .A1(n35355), .B0(n35368), .B1(n35354), .Y(
        n35356) );
  OR2XL U37130 ( .A(n35549), .B(n35356), .Y(n16277) );
  AOI2BB1XL U37131 ( .A0N(n35365), .A1N(n35358), .B0(n35357), .Y(n35359) );
  OAI2BB2XL U37132 ( .B0(conv_1[188]), .B1(n35359), .A0N(conv_1[188]), .A1N(
        n35359), .Y(n35361) );
  INVXL U37133 ( .A(conv_1[188]), .Y(n35360) );
  OAI22XL U37134 ( .A0(n36009), .A1(n35361), .B0(n35368), .B1(n35360), .Y(
        n35362) );
  OR2XL U37135 ( .A(n35549), .B(n35362), .Y(n16275) );
  OAI2BB2XL U37136 ( .B0(conv_1[190]), .B1(n35366), .A0N(conv_1[190]), .A1N(
        n35366), .Y(n35369) );
  OAI22XL U37137 ( .A0(n36009), .A1(n35369), .B0(n35368), .B1(n35367), .Y(
        n35370) );
  OR2XL U37138 ( .A(n35549), .B(n35370), .Y(n16273) );
  AOI2BB1XL U37139 ( .A0N(n35379), .A1N(n35372), .B0(n35371), .Y(n35373) );
  OAI2BB2XL U37140 ( .B0(conv_1[203]), .B1(n35373), .A0N(conv_1[203]), .A1N(
        n35373), .Y(n35375) );
  OAI2BB2XL U37141 ( .B0(n16654), .B1(n35375), .A0N(n35374), .A1N(conv_1[203]), 
        .Y(n35376) );
  OR2XL U37142 ( .A(n35549), .B(n35376), .Y(n16260) );
  AOI2BB1XL U37143 ( .A0N(n35379), .A1N(n35378), .B0(n35377), .Y(n35380) );
  OAI2BB2XL U37144 ( .B0(conv_1[205]), .B1(n35380), .A0N(conv_1[205]), .A1N(
        n35380), .Y(n35382) );
  OAI22XL U37145 ( .A0(n36009), .A1(n35382), .B0(n35384), .B1(n35381), .Y(
        n35383) );
  OR2XL U37146 ( .A(n35549), .B(n35383), .Y(n16258) );
  AOI32XL U37147 ( .A0(n35385), .A1(n35384), .A2(n35386), .B0(n36009), .B1(
        n35384), .Y(n35389) );
  AOI31XL U37148 ( .A0(n34028), .A1(n35387), .A2(n35386), .B0(n35549), .Y(
        n35388) );
  OAI2BB1XL U37149 ( .A0N(conv_1[206]), .A1N(n35389), .B0(n35388), .Y(n16257)
         );
  AOI2BB1XL U37150 ( .A0N(n35392), .A1N(n35391), .B0(n35390), .Y(n35393) );
  OAI2BB2XL U37151 ( .B0(conv_1[217]), .B1(n35393), .A0N(conv_1[217]), .A1N(
        n35393), .Y(n35396) );
  OAI22XL U37152 ( .A0(n36009), .A1(n35396), .B0(n35395), .B1(n35394), .Y(
        n35397) );
  OR2XL U37153 ( .A(n35549), .B(n35397), .Y(n16246) );
  AOI32XL U37154 ( .A0(n35399), .A1(n35408), .A2(n35398), .B0(n36001), .B1(
        n35408), .Y(n35402) );
  AOI31XL U37155 ( .A0(n32181), .A1(n35400), .A2(n35399), .B0(n35549), .Y(
        n35401) );
  OAI2BB1XL U37156 ( .A0N(conv_1[232]), .A1N(n35402), .B0(n35401), .Y(n16231)
         );
  AOI21XL U37157 ( .A0(n35405), .A1(n35404), .B0(n35403), .Y(n35406) );
  OAI2BB2XL U37158 ( .B0(conv_1[234]), .B1(n35406), .A0N(conv_1[234]), .A1N(
        n35406), .Y(n35409) );
  OAI22XL U37159 ( .A0(n36042), .A1(n35409), .B0(n35408), .B1(n35407), .Y(
        n35410) );
  OR2XL U37160 ( .A(n35549), .B(n35410), .Y(n16229) );
  NAND2XL U37161 ( .A(conv_1[249]), .B(n35411), .Y(n35413) );
  AOI21XL U37162 ( .A0(n35414), .A1(n35413), .B0(n35412), .Y(n35415) );
  OAI2BB2XL U37163 ( .B0(conv_1[250]), .B1(n35415), .A0N(conv_1[250]), .A1N(
        n35415), .Y(n35418) );
  OAI22XL U37164 ( .A0(n35419), .A1(n35418), .B0(n35417), .B1(n35416), .Y(
        n35420) );
  OR2XL U37165 ( .A(n35549), .B(n35420), .Y(n16213) );
  AOI32XL U37166 ( .A0(n35422), .A1(n35426), .A2(n35421), .B0(n36009), .B1(
        n35426), .Y(n35425) );
  AOI31XL U37167 ( .A0(n36020), .A1(n35423), .A2(n35422), .B0(n35549), .Y(
        n35424) );
  OAI2BB1XL U37168 ( .A0N(conv_1[278]), .A1N(n35425), .B0(n35424), .Y(n16185)
         );
  AOI32XL U37169 ( .A0(n35427), .A1(n35426), .A2(n35428), .B0(n16655), .B1(
        n35426), .Y(n35431) );
  OAI2BB1XL U37170 ( .A0N(conv_1[281]), .A1N(n35431), .B0(n35430), .Y(n16182)
         );
  AOI2BB1XL U37171 ( .A0N(n35434), .A1N(n35433), .B0(n35432), .Y(n35435) );
  OAI2BB2XL U37172 ( .B0(conv_1[338]), .B1(n35435), .A0N(conv_1[338]), .A1N(
        n35435), .Y(n35438) );
  OAI22XL U37173 ( .A0(n36001), .A1(n35438), .B0(n35437), .B1(n35436), .Y(
        n35439) );
  OR2XL U37174 ( .A(n35549), .B(n35439), .Y(n16125) );
  AOI21XL U37175 ( .A0(n35442), .A1(n35441), .B0(n35440), .Y(n35443) );
  OAI2BB2XL U37176 ( .B0(conv_1[354]), .B1(n35443), .A0N(conv_1[354]), .A1N(
        n35443), .Y(n35445) );
  OAI22XL U37177 ( .A0(n34389), .A1(n35445), .B0(n35447), .B1(n35444), .Y(
        n35446) );
  OR2XL U37178 ( .A(n35549), .B(n35446), .Y(n16109) );
  AOI32XL U37179 ( .A0(n35448), .A1(n35447), .A2(n35449), .B0(n36042), .B1(
        n35447), .Y(n35452) );
  AOI31XL U37180 ( .A0(n33778), .A1(n35450), .A2(n35449), .B0(n35549), .Y(
        n35451) );
  OAI2BB1XL U37181 ( .A0N(conv_1[356]), .A1N(n35452), .B0(n35451), .Y(n16107)
         );
  AOI2BB1XL U37182 ( .A0N(n35455), .A1N(n35454), .B0(n35453), .Y(n35456) );
  OAI2BB2XL U37183 ( .B0(conv_1[368]), .B1(n35456), .A0N(conv_1[368]), .A1N(
        n35456), .Y(n35459) );
  OAI22XL U37184 ( .A0(n36001), .A1(n35459), .B0(n35458), .B1(n35457), .Y(
        n35460) );
  OR2XL U37185 ( .A(n35549), .B(n35460), .Y(n16095) );
  AOI2BB1XL U37186 ( .A0N(n35463), .A1N(n35462), .B0(n35461), .Y(n35464) );
  OAI2BB2XL U37187 ( .B0(conv_1[383]), .B1(n35464), .A0N(conv_1[383]), .A1N(
        n35464), .Y(n35467) );
  OAI22XL U37188 ( .A0(n36001), .A1(n35467), .B0(n35466), .B1(n35465), .Y(
        n35468) );
  OR2XL U37189 ( .A(n35549), .B(n35468), .Y(n16080) );
  AOI21XL U37190 ( .A0(n35471), .A1(n35470), .B0(n35469), .Y(n35472) );
  OAI2BB2XL U37191 ( .B0(conv_1[399]), .B1(n35472), .A0N(conv_1[399]), .A1N(
        n35472), .Y(n35474) );
  OAI22XL U37192 ( .A0(n36001), .A1(n35474), .B0(n35477), .B1(n35473), .Y(
        n35475) );
  OR2XL U37193 ( .A(n35549), .B(n35475), .Y(n16064) );
  INVXL U37194 ( .A(n35476), .Y(n35478) );
  AOI32XL U37195 ( .A0(n35478), .A1(n35477), .A2(n35479), .B0(n16655), .B1(
        n35477), .Y(n35482) );
  OAI2BB1XL U37196 ( .A0N(conv_1[401]), .A1N(n35482), .B0(n35481), .Y(n16062)
         );
  XOR2XL U37197 ( .A(n35484), .B(n35483), .Y(n35485) );
  OAI2BB2XL U37198 ( .B0(conv_1[409]), .B1(n35485), .A0N(conv_1[409]), .A1N(
        n35485), .Y(n35488) );
  OAI22XL U37199 ( .A0(n16654), .A1(n35488), .B0(n35487), .B1(n35486), .Y(
        n35490) );
  NAND2BXL U37200 ( .AN(n35490), .B(n35489), .Y(n16054) );
  AOI2BB1XL U37201 ( .A0N(n35493), .A1N(n35492), .B0(n35491), .Y(n35494) );
  OAI2BB2XL U37202 ( .B0(conv_1[412]), .B1(n35494), .A0N(conv_1[412]), .A1N(
        n35494), .Y(n35496) );
  OAI2BB2XL U37203 ( .B0(n16654), .B1(n35496), .A0N(n35495), .A1N(conv_1[412]), 
        .Y(n35497) );
  OR2XL U37204 ( .A(n35549), .B(n35497), .Y(n16051) );
  AOI21XL U37205 ( .A0(intadd_1_n1), .A1(intadd_1_B_2_), .B0(n35501), .Y(
        n35502) );
  OAI2BB2XL U37206 ( .B0(conv_1[426]), .B1(n35502), .A0N(conv_1[426]), .A1N(
        n35502), .Y(n35505) );
  OAI22XL U37207 ( .A0(n36001), .A1(n35505), .B0(n35504), .B1(n35503), .Y(
        n35506) );
  OR2XL U37208 ( .A(n35549), .B(n35506), .Y(n16037) );
  AOI2BB1XL U37209 ( .A0N(intadd_1_B_2_), .A1N(n35508), .B0(n35507), .Y(n35509) );
  OAI2BB2XL U37210 ( .B0(conv_1[431]), .B1(n35509), .A0N(conv_1[431]), .A1N(
        n35509), .Y(n35511) );
  OAI2BB2XL U37211 ( .B0(n36009), .B1(n35511), .A0N(n35510), .A1N(conv_1[431]), 
        .Y(n35512) );
  OR2XL U37212 ( .A(n35549), .B(n35512), .Y(n16032) );
  AOI2BB1XL U37213 ( .A0N(n35515), .A1N(n35514), .B0(n35513), .Y(n35516) );
  OAI2BB2XL U37214 ( .B0(conv_1[445]), .B1(n35516), .A0N(conv_1[445]), .A1N(
        n35516), .Y(n35518) );
  OAI2BB2XL U37215 ( .B0(n16654), .B1(n35518), .A0N(n35517), .A1N(conv_1[445]), 
        .Y(n35519) );
  OR2XL U37216 ( .A(n35549), .B(n35519), .Y(n16018) );
  AOI32XL U37217 ( .A0(n35521), .A1(n35520), .A2(n35522), .B0(n16655), .B1(
        n35520), .Y(n35525) );
  AOI31XL U37218 ( .A0(n36020), .A1(n35523), .A2(n35522), .B0(n35549), .Y(
        n35524) );
  OAI2BB1XL U37219 ( .A0N(conv_1[446]), .A1N(n35525), .B0(n35524), .Y(n16017)
         );
  AOI2BB1XL U37220 ( .A0N(n35541), .A1N(n35527), .B0(n35526), .Y(n35528) );
  OAI2BB2XL U37221 ( .B0(conv_1[486]), .B1(n35528), .A0N(conv_1[486]), .A1N(
        n35528), .Y(n35530) );
  OAI22XL U37222 ( .A0(n16654), .A1(n35530), .B0(n35544), .B1(n35529), .Y(
        n35531) );
  OR2XL U37223 ( .A(n35549), .B(n35531), .Y(n15977) );
  AOI21XL U37224 ( .A0(n35534), .A1(n35533), .B0(n35532), .Y(n35535) );
  OAI2BB2XL U37225 ( .B0(conv_1[487]), .B1(n35535), .A0N(conv_1[487]), .A1N(
        n35535), .Y(n35537) );
  OAI22XL U37226 ( .A0(n16654), .A1(n35537), .B0(n35544), .B1(n35536), .Y(
        n35538) );
  OR2XL U37227 ( .A(n35549), .B(n35538), .Y(n15976) );
  AOI2BB1XL U37228 ( .A0N(n35541), .A1N(n35540), .B0(n35539), .Y(n35542) );
  OAI2BB2XL U37229 ( .B0(conv_1[488]), .B1(n35542), .A0N(conv_1[488]), .A1N(
        n35542), .Y(n35545) );
  INVXL U37230 ( .A(conv_1[488]), .Y(n35543) );
  OAI22XL U37231 ( .A0(n36001), .A1(n35545), .B0(n35544), .B1(n35543), .Y(
        n35546) );
  OR2XL U37232 ( .A(n35549), .B(n35546), .Y(n15975) );
  AOI32XL U37233 ( .A0(n35548), .A1(n35547), .A2(n35550), .B0(n16654), .B1(
        n35547), .Y(n35553) );
  AOI31XL U37234 ( .A0(n33778), .A1(n35551), .A2(n35550), .B0(n35549), .Y(
        n35552) );
  OAI2BB1XL U37235 ( .A0N(conv_1[521]), .A1N(n35553), .B0(n35552), .Y(n15942)
         );
  INVXL U37236 ( .A(n35554), .Y(n35555) );
  AOI32XL U37237 ( .A0(n35557), .A1(n35630), .A2(n35555), .B0(n36001), .B1(
        n35630), .Y(n35560) );
  INVXL U37238 ( .A(n35566), .Y(n35556) );
  AOI31XL U37239 ( .A0(n32181), .A1(n35558), .A2(n35557), .B0(n35556), .Y(
        n35559) );
  OAI2BB1XL U37240 ( .A0N(conv_3[167]), .A1N(n35560), .B0(n35559), .Y(n15840)
         );
  AOI32XL U37241 ( .A0(n35562), .A1(n35743), .A2(n35561), .B0(n36001), .B1(
        n35743), .Y(n35568) );
  OAI31XL U37242 ( .A0(n35565), .A1(n35564), .A2(n16654), .B0(n35563), .Y(
        n35567) );
  OAI2BB1XL U37243 ( .A0N(n35568), .A1N(n35567), .B0(n35566), .Y(n15830) );
  XOR2XL U37244 ( .A(n35570), .B(n35569), .Y(n35571) );
  OAI2BB2XL U37245 ( .B0(conv_3[123]), .B1(n35571), .A0N(conv_3[123]), .A1N(
        n35571), .Y(n35573) );
  OAI2BB2XL U37246 ( .B0(n16654), .B1(n35573), .A0N(n35572), .A1N(conv_3[123]), 
        .Y(n35575) );
  NAND2BXL U37247 ( .AN(n35575), .B(n35574), .Y(n15807) );
  AOI32XL U37248 ( .A0(n35577), .A1(n35576), .A2(n35578), .B0(n16655), .B1(
        n35576), .Y(n35581) );
  AOI31XL U37249 ( .A0(n36020), .A1(n35579), .A2(n35578), .B0(n16653), .Y(
        n35580) );
  OAI2BB1XL U37250 ( .A0N(conv_3[26]), .A1N(n35581), .B0(n35580), .Y(n15727)
         );
  INVXL U37251 ( .A(n35582), .Y(n35583) );
  AOI32XL U37252 ( .A0(n35584), .A1(n35594), .A2(n35583), .B0(n36009), .B1(
        n35594), .Y(n35587) );
  AOI31XL U37253 ( .A0(n36020), .A1(n35585), .A2(n35584), .B0(n16653), .Y(
        n35586) );
  OAI2BB1XL U37254 ( .A0N(conv_3[35]), .A1N(n35587), .B0(n35586), .Y(n15723)
         );
  AOI21XL U37255 ( .A0(n35591), .A1(n35590), .B0(n35589), .Y(n35592) );
  OAI2BB2XL U37256 ( .B0(conv_3[38]), .B1(n35592), .A0N(conv_3[38]), .A1N(
        n35592), .Y(n35595) );
  OAI22XL U37257 ( .A0(n36009), .A1(n35595), .B0(n35594), .B1(n35593), .Y(
        n35596) );
  OR2XL U37258 ( .A(n16653), .B(n35596), .Y(n15720) );
  NAND2XL U37259 ( .A(n35599), .B(n35600), .Y(n35597) );
  AOI32XL U37260 ( .A0(n35601), .A1(n35598), .A2(n35597), .B0(n36009), .B1(
        n35598), .Y(n35604) );
  AOI21XL U37261 ( .A0(n35600), .A1(n35599), .B0(conv_3[67]), .Y(n35602) );
  AOI31XL U37262 ( .A0(n31735), .A1(n35602), .A2(n35601), .B0(n16653), .Y(
        n35603) );
  OAI2BB1XL U37263 ( .A0N(conv_3[67]), .A1N(n35604), .B0(n35603), .Y(n15701)
         );
  AOI21XL U37264 ( .A0(n35607), .A1(n35606), .B0(n35605), .Y(n35608) );
  OAI2BB2XL U37265 ( .B0(conv_3[84]), .B1(n35608), .A0N(conv_3[84]), .A1N(
        n35608), .Y(n35611) );
  OAI22XL U37266 ( .A0(n34389), .A1(n35611), .B0(n35610), .B1(n35609), .Y(
        n35612) );
  OR2XL U37267 ( .A(n16653), .B(n35612), .Y(n15689) );
  AOI21XL U37268 ( .A0(n35615), .A1(n35614), .B0(n35613), .Y(n35616) );
  OAI2BB2XL U37269 ( .B0(conv_3[99]), .B1(n35616), .A0N(conv_3[99]), .A1N(
        n35616), .Y(n35619) );
  OAI22XL U37270 ( .A0(n36042), .A1(n35619), .B0(n35618), .B1(n35617), .Y(
        n35620) );
  OR2XL U37271 ( .A(n31384), .B(n35620), .Y(n15679) );
  AOI21XL U37272 ( .A0(n35623), .A1(n35622), .B0(n35621), .Y(n35624) );
  OAI2BB2XL U37273 ( .B0(conv_3[127]), .B1(n35624), .A0N(conv_3[127]), .A1N(
        n35624), .Y(n35627) );
  OAI22XL U37274 ( .A0(n36009), .A1(n35627), .B0(n35626), .B1(n35625), .Y(
        n35628) );
  OR2XL U37275 ( .A(n16653), .B(n35628), .Y(n15661) );
  AOI32XL U37276 ( .A0(n35631), .A1(n35630), .A2(n35629), .B0(n36042), .B1(
        n35630), .Y(n35634) );
  AOI2BB1XL U37277 ( .A0N(n35639), .A1N(n35638), .B0(n35637), .Y(n35640) );
  OAI2BB2XL U37278 ( .B0(conv_3[175]), .B1(n35640), .A0N(conv_3[175]), .A1N(
        n35640), .Y(n35642) );
  OAI2BB2XL U37279 ( .B0(n36001), .B1(n35642), .A0N(n35641), .A1N(conv_3[175]), 
        .Y(n35643) );
  OR2XL U37280 ( .A(n16653), .B(n35643), .Y(n15628) );
  INVXL U37281 ( .A(n35644), .Y(n35645) );
  AOI32XL U37282 ( .A0(n35647), .A1(n35646), .A2(n35645), .B0(n36001), .B1(
        n35646), .Y(n35650) );
  AOI2BB1XL U37283 ( .A0N(n35653), .A1N(n35652), .B0(n35651), .Y(n35654) );
  OAI2BB2XL U37284 ( .B0(conv_3[205]), .B1(n35654), .A0N(conv_3[205]), .A1N(
        n35654), .Y(n35656) );
  OAI2BB2XL U37285 ( .B0(n34389), .B1(n35656), .A0N(n35655), .A1N(conv_3[205]), 
        .Y(n35657) );
  OR2XL U37286 ( .A(n31384), .B(n35657), .Y(n15608) );
  AOI2BB1XL U37287 ( .A0N(n35660), .A1N(n35659), .B0(n35658), .Y(n35661) );
  OAI2BB2XL U37288 ( .B0(conv_3[216]), .B1(n35661), .A0N(conv_3[216]), .A1N(
        n35661), .Y(n35663) );
  OAI2BB2XL U37289 ( .B0(n16658), .B1(n35663), .A0N(n35662), .A1N(conv_3[216]), 
        .Y(n35664) );
  OR2XL U37290 ( .A(n16653), .B(n35664), .Y(n15602) );
  AOI32XL U37291 ( .A0(n35666), .A1(n35665), .A2(n35667), .B0(n34389), .B1(
        n35665), .Y(n35670) );
  AOI2BB1XL U37292 ( .A0N(n35673), .A1N(n35672), .B0(n35671), .Y(n35674) );
  OAI2BB2XL U37293 ( .B0(conv_3[233]), .B1(n35674), .A0N(conv_3[233]), .A1N(
        n35674), .Y(n35677) );
  OAI22XL U37294 ( .A0(n36001), .A1(n35677), .B0(n35676), .B1(n35675), .Y(
        n35678) );
  OR2XL U37295 ( .A(n16653), .B(n35678), .Y(n15590) );
  AOI2BB1XL U37296 ( .A0N(n35693), .A1N(n35680), .B0(n35679), .Y(n35681) );
  OAI2BB2XL U37297 ( .B0(conv_3[246]), .B1(n35681), .A0N(conv_3[246]), .A1N(
        n35681), .Y(n35683) );
  OAI22XL U37298 ( .A0(n36001), .A1(n35683), .B0(n35706), .B1(n35682), .Y(
        n35684) );
  OR2XL U37299 ( .A(n16653), .B(n35684), .Y(n15582) );
  AOI21XL U37300 ( .A0(n35700), .A1(n35686), .B0(n35685), .Y(n35687) );
  OAI2BB2XL U37301 ( .B0(conv_3[247]), .B1(n35687), .A0N(conv_3[247]), .A1N(
        n35687), .Y(n35689) );
  OAI22XL U37302 ( .A0(n36001), .A1(n35689), .B0(n35706), .B1(n35688), .Y(
        n35690) );
  OR2XL U37303 ( .A(n31384), .B(n35690), .Y(n15581) );
  AOI2BB1XL U37304 ( .A0N(n35693), .A1N(n35692), .B0(n35691), .Y(n35694) );
  OAI2BB2XL U37305 ( .B0(conv_3[248]), .B1(n35694), .A0N(conv_3[248]), .A1N(
        n35694), .Y(n35696) );
  OAI22XL U37306 ( .A0(n36001), .A1(n35696), .B0(n35706), .B1(n35695), .Y(
        n35697) );
  OR2XL U37307 ( .A(n16653), .B(n35697), .Y(n15580) );
  AOI21XL U37308 ( .A0(n35700), .A1(n35699), .B0(n35698), .Y(n35701) );
  OAI2BB2XL U37309 ( .B0(conv_3[249]), .B1(n35701), .A0N(conv_3[249]), .A1N(
        n35701), .Y(n35703) );
  OAI22XL U37310 ( .A0(n36001), .A1(n35703), .B0(n35706), .B1(n35702), .Y(
        n35704) );
  OR2XL U37311 ( .A(n16653), .B(n35704), .Y(n15579) );
  INVXL U37312 ( .A(n35705), .Y(n35707) );
  AOI32XL U37313 ( .A0(n35707), .A1(n35706), .A2(n35708), .B0(n36009), .B1(
        n35706), .Y(n35711) );
  OAI2BB1XL U37314 ( .A0N(conv_3[251]), .A1N(n35711), .B0(n35710), .Y(n15577)
         );
  AOI32XL U37315 ( .A0(n35714), .A1(n35713), .A2(n35712), .B0(n16654), .B1(
        n35713), .Y(n35717) );
  AOI31XL U37316 ( .A0(n32611), .A1(n35715), .A2(n35714), .B0(n16653), .Y(
        n35716) );
  OAI2BB1XL U37317 ( .A0N(conv_3[265]), .A1N(n35717), .B0(n35716), .Y(n15568)
         );
  AOI2BB1XL U37318 ( .A0N(n35720), .A1N(n35719), .B0(n35718), .Y(n35721) );
  OAI2BB2XL U37319 ( .B0(conv_3[293]), .B1(n35721), .A0N(conv_3[293]), .A1N(
        n35721), .Y(n35723) );
  OAI22XL U37320 ( .A0(n36001), .A1(n35723), .B0(n35726), .B1(n35722), .Y(
        n35724) );
  OR2XL U37321 ( .A(n16653), .B(n35724), .Y(n15550) );
  AOI32XL U37322 ( .A0(n35727), .A1(n35726), .A2(n35725), .B0(n36009), .B1(
        n35726), .Y(n35730) );
  OAI2BB1XL U37323 ( .A0N(conv_3[294]), .A1N(n35730), .B0(n35729), .Y(n15549)
         );
  AOI21XL U37324 ( .A0(n35733), .A1(n35732), .B0(n35731), .Y(n35734) );
  OAI2BB2XL U37325 ( .B0(conv_3[307]), .B1(n35734), .A0N(conv_3[307]), .A1N(
        n35734), .Y(n35737) );
  OAI22XL U37326 ( .A0(n16654), .A1(n35737), .B0(n35736), .B1(n35735), .Y(
        n35738) );
  OR2XL U37327 ( .A(n31384), .B(n35738), .Y(n15541) );
  OAI2BB2XL U37328 ( .B0(conv_3[323]), .B1(n35741), .A0N(conv_3[323]), .A1N(
        n35741), .Y(n35744) );
  OAI22XL U37329 ( .A0(n36001), .A1(n35744), .B0(n35743), .B1(n35742), .Y(
        n35745) );
  OR2XL U37330 ( .A(n16653), .B(n35745), .Y(n15530) );
  INVXL U37331 ( .A(n35746), .Y(n35747) );
  AOI32XL U37332 ( .A0(n35749), .A1(n35748), .A2(n35747), .B0(n36001), .B1(
        n35748), .Y(n35752) );
  AOI31XL U37333 ( .A0(n36020), .A1(n35750), .A2(n35749), .B0(n16653), .Y(
        n35751) );
  OAI2BB1XL U37334 ( .A0N(conv_3[335]), .A1N(n35752), .B0(n35751), .Y(n15523)
         );
  OAI2BB2XL U37335 ( .B0(conv_3[336]), .B1(n35755), .A0N(conv_3[336]), .A1N(
        n35755), .Y(n35757) );
  OAI2BB2XL U37336 ( .B0(n16654), .B1(n35757), .A0N(n35756), .A1N(conv_3[336]), 
        .Y(n35758) );
  OR2XL U37337 ( .A(n16653), .B(n35758), .Y(n15522) );
  AOI21XL U37338 ( .A0(n35761), .A1(n35760), .B0(n35759), .Y(n35762) );
  OAI2BB2XL U37339 ( .B0(conv_3[369]), .B1(n35762), .A0N(conv_3[369]), .A1N(
        n35762), .Y(n35765) );
  OAI22XL U37340 ( .A0(n16654), .A1(n35765), .B0(n35764), .B1(n35763), .Y(
        n35766) );
  OR2XL U37341 ( .A(n16653), .B(n35766), .Y(n15499) );
  AOI21XL U37342 ( .A0(n35775), .A1(n35768), .B0(n35767), .Y(n35769) );
  OAI2BB2XL U37343 ( .B0(conv_3[427]), .B1(n35769), .A0N(conv_3[427]), .A1N(
        n35769), .Y(n35771) );
  OAI22XL U37344 ( .A0(n36042), .A1(n35771), .B0(n35778), .B1(n35770), .Y(
        n35772) );
  OR2XL U37345 ( .A(n16653), .B(n35772), .Y(n15461) );
  AOI21XL U37346 ( .A0(n35775), .A1(n35774), .B0(n35773), .Y(n35776) );
  OAI2BB2XL U37347 ( .B0(conv_3[429]), .B1(n35776), .A0N(conv_3[429]), .A1N(
        n35776), .Y(n35779) );
  OAI22XL U37348 ( .A0(n36042), .A1(n35779), .B0(n35778), .B1(n35777), .Y(
        n35780) );
  OR2XL U37349 ( .A(n16653), .B(n35780), .Y(n15459) );
  AOI21XL U37350 ( .A0(n35789), .A1(n35782), .B0(n35781), .Y(n35783) );
  OAI2BB2XL U37351 ( .B0(conv_3[442]), .B1(n35783), .A0N(conv_3[442]), .A1N(
        n35783), .Y(n35785) );
  OAI22XL U37352 ( .A0(n36042), .A1(n35785), .B0(n35792), .B1(n35784), .Y(
        n35786) );
  OR2XL U37353 ( .A(n16653), .B(n35786), .Y(n15451) );
  AOI21XL U37354 ( .A0(n35789), .A1(n35788), .B0(n35787), .Y(n35790) );
  OAI2BB2XL U37355 ( .B0(conv_3[444]), .B1(n35790), .A0N(conv_3[444]), .A1N(
        n35790), .Y(n35793) );
  OAI22XL U37356 ( .A0(n36042), .A1(n35793), .B0(n35792), .B1(n35791), .Y(
        n35794) );
  OR2XL U37357 ( .A(n16653), .B(n35794), .Y(n15449) );
  INVXL U37358 ( .A(n35795), .Y(n35796) );
  OAI221XL U37359 ( .A0(n35797), .A1(n16658), .B0(n35796), .B1(n16655), .C0(
        n35805), .Y(n35800) );
  AOI31XL U37360 ( .A0(n36020), .A1(n35798), .A2(n35797), .B0(n16653), .Y(
        n35799) );
  OAI2BB1XL U37361 ( .A0N(n35800), .A1N(conv_3[455]), .B0(n35799), .Y(n15443)
         );
  OAI2BB2XL U37362 ( .B0(conv_3[458]), .B1(n35803), .A0N(conv_3[458]), .A1N(
        n35803), .Y(n35806) );
  OAI22XL U37363 ( .A0(n36042), .A1(n35806), .B0(n35805), .B1(n35804), .Y(
        n35807) );
  OR2XL U37364 ( .A(n16653), .B(n35807), .Y(n15440) );
  AOI2BB1XL U37365 ( .A0N(n35810), .A1N(n35809), .B0(n35808), .Y(n35811) );
  OAI2BB2XL U37366 ( .B0(conv_3[471]), .B1(n35811), .A0N(conv_3[471]), .A1N(
        n35811), .Y(n35814) );
  OAI22XL U37367 ( .A0(n16655), .A1(n35814), .B0(n35813), .B1(n35812), .Y(
        n35815) );
  OR2XL U37368 ( .A(n16653), .B(n35815), .Y(n15432) );
  NAND2XL U37369 ( .A(n35831), .B(n35822), .Y(n35816) );
  AOI32XL U37370 ( .A0(n35816), .A1(n35826), .A2(n35817), .B0(n16658), .B1(
        n35826), .Y(n35820) );
  AOI21XL U37371 ( .A0(n35831), .A1(n35822), .B0(conv_3[486]), .Y(n35818) );
  AOI31XL U37372 ( .A0(n24378), .A1(n35818), .A2(n35817), .B0(n16653), .Y(
        n35819) );
  OAI2BB1XL U37373 ( .A0N(conv_3[486]), .A1N(n35820), .B0(n35819), .Y(n15422)
         );
  OAI32XL U37374 ( .A0(n35823), .A1(conv_3[486]), .A2(n35822), .B0(n35831), 
        .B1(n35821), .Y(n35824) );
  OAI2BB2XL U37375 ( .B0(conv_3[487]), .B1(n35824), .A0N(conv_3[487]), .A1N(
        n35824), .Y(n35827) );
  OAI22XL U37376 ( .A0(n16655), .A1(n35827), .B0(n35826), .B1(n35825), .Y(
        n35828) );
  OR2XL U37377 ( .A(n16653), .B(n35828), .Y(n15421) );
  AOI2BB1XL U37378 ( .A0N(n35831), .A1N(n35830), .B0(n35829), .Y(n35832) );
  OAI2BB2XL U37379 ( .B0(conv_3[490]), .B1(n35832), .A0N(conv_3[490]), .A1N(
        n35832), .Y(n35834) );
  OAI2BB2XL U37380 ( .B0(n34389), .B1(n35834), .A0N(n35833), .A1N(conv_3[490]), 
        .Y(n35835) );
  OR2XL U37381 ( .A(n16653), .B(n35835), .Y(n15418) );
  AOI2BB1XL U37382 ( .A0N(n35838), .A1N(n35837), .B0(n35836), .Y(n35839) );
  OAI2BB2XL U37383 ( .B0(conv_3[501]), .B1(n35839), .A0N(conv_3[501]), .A1N(
        n35839), .Y(n35842) );
  OAI22XL U37384 ( .A0(n16655), .A1(n35842), .B0(n35841), .B1(n35840), .Y(
        n35843) );
  OR2XL U37385 ( .A(n16653), .B(n35843), .Y(n15412) );
  INVXL U37386 ( .A(n35844), .Y(n35845) );
  AOI32XL U37387 ( .A0(n35849), .A1(n35846), .A2(n35845), .B0(n16655), .B1(
        n35846), .Y(n35852) );
  INVXL U37388 ( .A(n35847), .Y(n35848) );
  AOI31XL U37389 ( .A0(n33982), .A1(n35850), .A2(n35849), .B0(n35848), .Y(
        n35851) );
  OAI2BB1XL U37390 ( .A0N(conv_2[61]), .A1N(n35852), .B0(n35851), .Y(n15343)
         );
  OAI2BB2XL U37391 ( .B0(n18913), .B1(n35855), .A0N(n35854), .A1N(conv_2[1]), 
        .Y(intadd_0_CI) );
  AOI21XL U37392 ( .A0(n35862), .A1(n35861), .B0(n35860), .Y(n35863) );
  OAI2BB2XL U37393 ( .B0(conv_2[39]), .B1(n35863), .A0N(conv_2[39]), .A1N(
        n35863), .Y(n35866) );
  OAI22XL U37394 ( .A0(n16654), .A1(n35866), .B0(n35865), .B1(n35864), .Y(
        n35867) );
  OR2XL U37395 ( .A(n16651), .B(n35867), .Y(n15179) );
  AOI2BB1XL U37396 ( .A0N(n35876), .A1N(n35869), .B0(n35868), .Y(n35870) );
  OAI2BB2XL U37397 ( .B0(conv_2[81]), .B1(n35870), .A0N(conv_2[81]), .A1N(
        n35870), .Y(n35872) );
  OAI22XL U37398 ( .A0(n36009), .A1(n35872), .B0(n35879), .B1(n35871), .Y(
        n35873) );
  OR2XL U37399 ( .A(n16651), .B(n35873), .Y(n15152) );
  AOI2BB1XL U37400 ( .A0N(n35876), .A1N(n35875), .B0(n35874), .Y(n35877) );
  OAI2BB2XL U37401 ( .B0(conv_2[83]), .B1(n35877), .A0N(conv_2[83]), .A1N(
        n35877), .Y(n35880) );
  OAI22XL U37402 ( .A0(n36042), .A1(n35880), .B0(n35879), .B1(n35878), .Y(
        n35881) );
  OR2XL U37403 ( .A(n16651), .B(n35881), .Y(n15150) );
  AOI21XL U37404 ( .A0(n35884), .A1(n35883), .B0(n35882), .Y(n35885) );
  OAI2BB2XL U37405 ( .B0(conv_2[112]), .B1(n35885), .A0N(conv_2[112]), .A1N(
        n35885), .Y(n35887) );
  OAI22XL U37406 ( .A0(n36001), .A1(n35887), .B0(n35894), .B1(n35886), .Y(
        n35888) );
  OR2XL U37407 ( .A(n16651), .B(n35888), .Y(n15131) );
  AOI2BB1XL U37408 ( .A0N(n35891), .A1N(n35890), .B0(n35889), .Y(n35892) );
  OAI2BB2XL U37409 ( .B0(conv_2[113]), .B1(n35892), .A0N(conv_2[113]), .A1N(
        n35892), .Y(n35895) );
  OAI22XL U37410 ( .A0(n36001), .A1(n35895), .B0(n35894), .B1(n35893), .Y(
        n35896) );
  OR2XL U37411 ( .A(n16651), .B(n35896), .Y(n15130) );
  AOI21XL U37412 ( .A0(n35899), .A1(n35898), .B0(n35897), .Y(n35900) );
  OAI2BB2XL U37413 ( .B0(conv_2[142]), .B1(n35900), .A0N(conv_2[142]), .A1N(
        n35900), .Y(n35903) );
  OAI22XL U37414 ( .A0(n34389), .A1(n35903), .B0(n35902), .B1(n35901), .Y(
        n35904) );
  OR2XL U37415 ( .A(n16651), .B(n35904), .Y(n15111) );
  AOI2BB1XL U37416 ( .A0N(n35907), .A1N(n35906), .B0(n35905), .Y(n35908) );
  OAI2BB2XL U37417 ( .B0(conv_2[143]), .B1(n35908), .A0N(conv_2[143]), .A1N(
        n35908), .Y(n35910) );
  OAI2BB2XL U37418 ( .B0(n16654), .B1(n35910), .A0N(n35909), .A1N(conv_2[143]), 
        .Y(n35911) );
  OR2XL U37419 ( .A(n16651), .B(n35911), .Y(n15110) );
  AOI2BB1XL U37420 ( .A0N(n35914), .A1N(n35913), .B0(n35912), .Y(n35915) );
  OAI2BB2XL U37421 ( .B0(conv_2[188]), .B1(n35915), .A0N(conv_2[188]), .A1N(
        n35915), .Y(n35918) );
  OAI22XL U37422 ( .A0(n36009), .A1(n35918), .B0(n35917), .B1(n35916), .Y(
        n35919) );
  OR2XL U37423 ( .A(n16651), .B(n35919), .Y(n15080) );
  AOI21XL U37424 ( .A0(n35928), .A1(n35921), .B0(n35920), .Y(n35922) );
  OAI2BB2XL U37425 ( .B0(conv_2[201]), .B1(n35922), .A0N(conv_2[201]), .A1N(
        n35922), .Y(n35924) );
  OAI22XL U37426 ( .A0(n36001), .A1(n35924), .B0(n35931), .B1(n35923), .Y(
        n35925) );
  OR2XL U37427 ( .A(n16651), .B(n35925), .Y(n15072) );
  AOI21XL U37428 ( .A0(n35928), .A1(n35927), .B0(n35926), .Y(n35929) );
  OAI2BB2XL U37429 ( .B0(conv_2[203]), .B1(n35929), .A0N(conv_2[203]), .A1N(
        n35929), .Y(n35932) );
  OAI22XL U37430 ( .A0(n36001), .A1(n35932), .B0(n35931), .B1(n35930), .Y(
        n35933) );
  OR2XL U37431 ( .A(n16651), .B(n35933), .Y(n15070) );
  AOI32XL U37432 ( .A0(n35935), .A1(n35934), .A2(n35936), .B0(n16658), .B1(
        n35934), .Y(n35939) );
  OAI2BB1XL U37433 ( .A0N(conv_2[221]), .A1N(n35939), .B0(n35938), .Y(n15057)
         );
  AOI2BB1XL U37434 ( .A0N(n35942), .A1N(n35941), .B0(n35940), .Y(n35943) );
  OAI2BB2XL U37435 ( .B0(conv_2[251]), .B1(n35943), .A0N(conv_2[251]), .A1N(
        n35943), .Y(n35946) );
  OAI22XL U37436 ( .A0(n36001), .A1(n35946), .B0(n35945), .B1(n35944), .Y(
        n35947) );
  OR2XL U37437 ( .A(n16651), .B(n35947), .Y(n15037) );
  AOI2BB1XL U37438 ( .A0N(n35950), .A1N(n35949), .B0(n35948), .Y(n35951) );
  OAI2BB2XL U37439 ( .B0(conv_2[280]), .B1(n35951), .A0N(conv_2[280]), .A1N(
        n35951), .Y(n35953) );
  OAI2BB2XL U37440 ( .B0(n16654), .B1(n35953), .A0N(n35952), .A1N(conv_2[280]), 
        .Y(n35954) );
  OR2XL U37441 ( .A(n16651), .B(n35954), .Y(n15018) );
  AOI2BB1XL U37442 ( .A0N(n35957), .A1N(n35956), .B0(n35955), .Y(n35958) );
  OAI2BB2XL U37443 ( .B0(conv_2[291]), .B1(n35958), .A0N(conv_2[291]), .A1N(
        n35958), .Y(n35960) );
  OAI2BB2XL U37444 ( .B0(n16654), .B1(n35960), .A0N(n35959), .A1N(conv_2[291]), 
        .Y(n35961) );
  OR2XL U37445 ( .A(n16651), .B(n35961), .Y(n15012) );
  AOI32XL U37446 ( .A0(n35964), .A1(n35963), .A2(n35962), .B0(n16654), .B1(
        n35963), .Y(n35967) );
  AOI31XL U37447 ( .A0(n33778), .A1(n35965), .A2(n35964), .B0(n16651), .Y(
        n35966) );
  OAI2BB1XL U37448 ( .A0N(conv_2[295]), .A1N(n35967), .B0(n35966), .Y(n15008)
         );
  AOI21XL U37449 ( .A0(n35970), .A1(n35969), .B0(n35968), .Y(n35971) );
  OAI2BB2XL U37450 ( .B0(conv_2[309]), .B1(n35971), .A0N(conv_2[309]), .A1N(
        n35971), .Y(n35973) );
  OAI22XL U37451 ( .A0(n16654), .A1(n35973), .B0(n35976), .B1(n35972), .Y(
        n35974) );
  OR2XL U37452 ( .A(n16651), .B(n35974), .Y(n14999) );
  AOI32XL U37453 ( .A0(n35977), .A1(n35976), .A2(n35975), .B0(n36042), .B1(
        n35976), .Y(n35980) );
  AOI31XL U37454 ( .A0(n36020), .A1(n35978), .A2(n35977), .B0(n16651), .Y(
        n35979) );
  OAI2BB1XL U37455 ( .A0N(conv_2[311]), .A1N(n35980), .B0(n35979), .Y(n14997)
         );
  AOI21XL U37456 ( .A0(n35983), .A1(n35982), .B0(n35981), .Y(n35984) );
  OAI2BB2XL U37457 ( .B0(conv_2[322]), .B1(n35984), .A0N(conv_2[322]), .A1N(
        n35984), .Y(n35987) );
  OAI22XL U37458 ( .A0(n36001), .A1(n35987), .B0(n35986), .B1(n35985), .Y(
        n35988) );
  OR2XL U37459 ( .A(n16651), .B(n35988), .Y(n14991) );
  AOI32XL U37460 ( .A0(n35990), .A1(n36003), .A2(n35989), .B0(n16654), .B1(
        n36003), .Y(n35993) );
  AOI31XL U37461 ( .A0(n36020), .A1(n35991), .A2(n35990), .B0(n16651), .Y(
        n35992) );
  OAI2BB1XL U37462 ( .A0N(conv_2[336]), .A1N(n35993), .B0(n35992), .Y(n14982)
         );
  OAI32XL U37463 ( .A0(n35997), .A1(conv_2[338]), .A2(n35996), .B0(n35995), 
        .B1(n35994), .Y(n35998) );
  OAI2BB2XL U37464 ( .B0(conv_2[339]), .B1(n35998), .A0N(conv_2[339]), .A1N(
        n35998), .Y(n36000) );
  OAI22XL U37465 ( .A0(n36001), .A1(n36000), .B0(n36003), .B1(n35999), .Y(
        n36002) );
  OR2XL U37466 ( .A(n16651), .B(n36002), .Y(n14979) );
  AOI32XL U37467 ( .A0(n36004), .A1(n36003), .A2(n36005), .B0(n16655), .B1(
        n36003), .Y(n36008) );
  AOI31XL U37468 ( .A0(n30090), .A1(n36006), .A2(n36005), .B0(n16651), .Y(
        n36007) );
  OAI2BB1XL U37469 ( .A0N(conv_2[341]), .A1N(n36008), .B0(n36007), .Y(n14977)
         );
  AOI32XL U37470 ( .A0(n36011), .A1(n36010), .A2(n36012), .B0(n36009), .B1(
        n36010), .Y(n36015) );
  AOI31XL U37471 ( .A0(n32656), .A1(n36013), .A2(n36012), .B0(n16651), .Y(
        n36014) );
  OAI2BB1XL U37472 ( .A0N(conv_2[356]), .A1N(n36015), .B0(n36014), .Y(n14967)
         );
  AOI32XL U37473 ( .A0(n36018), .A1(n36017), .A2(n36016), .B0(n34389), .B1(
        n36017), .Y(n36022) );
  AOI31XL U37474 ( .A0(n36020), .A1(n36019), .A2(n36018), .B0(n16651), .Y(
        n36021) );
  OAI2BB1XL U37475 ( .A0N(conv_2[366]), .A1N(n36022), .B0(n36021), .Y(n14962)
         );
  AOI21XL U37476 ( .A0(n36025), .A1(n36024), .B0(n36023), .Y(n36026) );
  OAI2BB2XL U37477 ( .B0(conv_2[382]), .B1(n36026), .A0N(conv_2[382]), .A1N(
        n36026), .Y(n36029) );
  OAI22XL U37478 ( .A0(n16654), .A1(n36029), .B0(n36028), .B1(n36027), .Y(
        n36030) );
  OR2XL U37479 ( .A(n16651), .B(n36030), .Y(n14951) );
  AOI32XL U37480 ( .A0(n36032), .A1(n36031), .A2(n36033), .B0(n36001), .B1(
        n36031), .Y(n36036) );
  AOI31XL U37481 ( .A0(n31735), .A1(n36034), .A2(n36033), .B0(n16651), .Y(
        n36035) );
  OAI2BB1XL U37482 ( .A0N(conv_2[401]), .A1N(n36036), .B0(n36035), .Y(n14937)
         );
  OAI2BB2XL U37483 ( .B0(conv_2[415]), .B1(n36039), .A0N(conv_2[415]), .A1N(
        n36039), .Y(n36041) );
  OAI22XL U37484 ( .A0(n36042), .A1(n36041), .B0(n36047), .B1(n36040), .Y(
        n36043) );
  OR2XL U37485 ( .A(n16651), .B(n36043), .Y(n14928) );
  OR2XL U37486 ( .A(n36045), .B(n36044), .Y(n36048) );
  NAND2XL U37487 ( .A(n36045), .B(n36044), .Y(n36046) );
  AOI32XL U37488 ( .A0(n36048), .A1(n36047), .A2(n36046), .B0(n16655), .B1(
        n36047), .Y(n36051) );
  OAI2BB1XL U37489 ( .A0N(conv_2[417]), .A1N(n36051), .B0(n36050), .Y(n14926)
         );
  AOI32XL U37490 ( .A0(n36054), .A1(n36053), .A2(n36052), .B0(n16654), .B1(
        n36053), .Y(n36058) );
  OAI2BB1XL U37491 ( .A0N(conv_2[429]), .A1N(n36058), .B0(n36057), .Y(n14919)
         );
  AOI2BB1XL U37492 ( .A0N(n36067), .A1N(n36060), .B0(n36059), .Y(n36061) );
  OAI2BB2XL U37493 ( .B0(conv_2[441]), .B1(n36061), .A0N(conv_2[441]), .A1N(
        n36061), .Y(n36063) );
  INVXL U37494 ( .A(conv_2[441]), .Y(n36062) );
  OAI22XL U37495 ( .A0(n34389), .A1(n36063), .B0(n36070), .B1(n36062), .Y(
        n36064) );
  AOI2BB1XL U37496 ( .A0N(n36067), .A1N(n36066), .B0(n36065), .Y(n36068) );
  OAI2BB2XL U37497 ( .B0(conv_2[443]), .B1(n36068), .A0N(conv_2[443]), .A1N(
        n36068), .Y(n36071) );
  INVXL U37498 ( .A(conv_2[443]), .Y(n36069) );
  OAI22XL U37499 ( .A0(n16655), .A1(n36071), .B0(n36070), .B1(n36069), .Y(
        n36072) );
  OR2XL U37500 ( .A(n16651), .B(n36072), .Y(n14910) );
  AOI2BB1XL U37501 ( .A0N(n36088), .A1N(n36074), .B0(n36073), .Y(n36075) );
  OAI2BB2XL U37502 ( .B0(conv_2[503]), .B1(n36075), .A0N(conv_2[503]), .A1N(
        n36075), .Y(n36077) );
  INVXL U37503 ( .A(conv_2[503]), .Y(n36076) );
  OAI22XL U37504 ( .A0(n34389), .A1(n36077), .B0(n36091), .B1(n36076), .Y(
        n36078) );
  AOI21XL U37505 ( .A0(n36081), .A1(n36080), .B0(n36079), .Y(n36082) );
  OAI2BB2XL U37506 ( .B0(conv_2[504]), .B1(n36082), .A0N(conv_2[504]), .A1N(
        n36082), .Y(n36084) );
  OAI22XL U37507 ( .A0(n16655), .A1(n36084), .B0(n36091), .B1(n36083), .Y(
        n36085) );
  OR2XL U37508 ( .A(n16651), .B(n36085), .Y(n14869) );
  AOI2BB1XL U37509 ( .A0N(n36088), .A1N(n36087), .B0(n36086), .Y(n36089) );
  OAI2BB2XL U37510 ( .B0(conv_2[505]), .B1(n36089), .A0N(conv_2[505]), .A1N(
        n36089), .Y(n36092) );
  OAI22XL U37511 ( .A0(n36001), .A1(n36092), .B0(n36091), .B1(n36090), .Y(
        n36093) );
  OR2XL U37512 ( .A(n16651), .B(n36093), .Y(n14868) );
  OAI2BB2XL U37513 ( .B0(n36136), .B1(n36124), .A0N(weight_2_bias_3[0]), .A1N(
        n36136), .Y(n14663) );
  INVXL U37514 ( .A(weight_2_bias_3[0]), .Y(n36125) );
  OAI2BB2XL U37515 ( .B0(n36136), .B1(n36125), .A0N(weight_2_bias_2[0]), .A1N(
        n36136), .Y(n14662) );
  INVXL U37516 ( .A(weight_2_bias_2[0]), .Y(n36126) );
  OAI2BB2XL U37517 ( .B0(n36126), .B1(n36136), .A0N(weight_2_bias_1[0]), .A1N(
        n36136), .Y(n14661) );
  OAI2BB2XL U37518 ( .B0(n36151), .B1(n36136), .A0N(weight_2_bias_3[5]), .A1N(
        n36136), .Y(n14660) );
  INVXL U37519 ( .A(weight_2_bias_3[5]), .Y(n36127) );
  OAI2BB2XL U37520 ( .B0(n36127), .B1(n36136), .A0N(weight_2_bias_2[5]), .A1N(
        n36136), .Y(n14659) );
  INVXL U37521 ( .A(weight_2_bias_2[5]), .Y(n36128) );
  OAI2BB2XL U37522 ( .B0(n36128), .B1(n36136), .A0N(weight_2_bias_1[5]), .A1N(
        n36136), .Y(n14658) );
  OAI2BB2XL U37523 ( .B0(n36148), .B1(n36136), .A0N(weight_2_bias_3[4]), .A1N(
        n36136), .Y(n14657) );
  INVXL U37524 ( .A(weight_2_bias_3[4]), .Y(n36129) );
  OAI2BB2XL U37525 ( .B0(n36129), .B1(n36136), .A0N(weight_2_bias_2[4]), .A1N(
        n36136), .Y(n14656) );
  INVXL U37526 ( .A(weight_2_bias_2[4]), .Y(n36130) );
  OAI2BB2XL U37527 ( .B0(n36130), .B1(n36136), .A0N(weight_2_bias_1[4]), .A1N(
        n36136), .Y(n14655) );
  OAI2BB2XL U37528 ( .B0(n36145), .B1(n36136), .A0N(weight_2_bias_3[3]), .A1N(
        n36136), .Y(n14654) );
  INVXL U37529 ( .A(weight_2_bias_3[3]), .Y(n36131) );
  OAI2BB2XL U37530 ( .B0(n36131), .B1(n36136), .A0N(weight_2_bias_2[3]), .A1N(
        n36136), .Y(n14653) );
  INVXL U37531 ( .A(weight_2_bias_2[3]), .Y(n36132) );
  OAI2BB2XL U37532 ( .B0(n36132), .B1(n36136), .A0N(weight_2_bias_1[3]), .A1N(
        n36136), .Y(n14652) );
  OAI2BB2XL U37533 ( .B0(n36142), .B1(n36136), .A0N(weight_2_bias_3[2]), .A1N(
        n36136), .Y(n14651) );
  INVXL U37534 ( .A(weight_2_bias_3[2]), .Y(n36133) );
  OAI2BB2XL U37535 ( .B0(n36133), .B1(n36136), .A0N(weight_2_bias_2[2]), .A1N(
        n36136), .Y(n14650) );
  INVXL U37536 ( .A(weight_2_bias_2[2]), .Y(n36134) );
  OAI2BB2XL U37537 ( .B0(n36134), .B1(n36136), .A0N(weight_2_bias_1[2]), .A1N(
        n36136), .Y(n14649) );
  OAI2BB2XL U37538 ( .B0(n36139), .B1(n36136), .A0N(weight_2_bias_3[1]), .A1N(
        n36136), .Y(n14648) );
  INVXL U37539 ( .A(weight_2_bias_3[1]), .Y(n36135) );
  OAI2BB2XL U37540 ( .B0(n36135), .B1(n36136), .A0N(weight_2_bias_2[1]), .A1N(
        n36136), .Y(n14647) );
  INVXL U37541 ( .A(weight_2_bias_2[1]), .Y(n36137) );
  OAI2BB2XL U37542 ( .B0(n36137), .B1(n36136), .A0N(weight_2_bias_1[1]), .A1N(
        n36136), .Y(n14646) );
  OAI2BB2XL U37543 ( .B0(n36153), .B1(n36138), .A0N(weight_1_bias_1[0]), .A1N(
        n36153), .Y(n14103) );
  OAI2BB2XL U37544 ( .B0(n36139), .B1(n36153), .A0N(weight_1_bias_3[1]), .A1N(
        n36153), .Y(n14102) );
  NAND2XL U37545 ( .A(weight_1_bias_2[1]), .B(n36153), .Y(n36140) );
  OAI2BB1XL U37546 ( .A0N(weight_1_bias_3[1]), .A1N(n36155), .B0(n36140), .Y(
        n14101) );
  NAND2XL U37547 ( .A(weight_1_bias_1[1]), .B(n36153), .Y(n36141) );
  OAI2BB1XL U37548 ( .A0N(weight_1_bias_2[1]), .A1N(n36155), .B0(n36141), .Y(
        n14100) );
  OAI2BB2XL U37549 ( .B0(n36142), .B1(n36153), .A0N(weight_1_bias_3[2]), .A1N(
        n36153), .Y(n14099) );
  NAND2XL U37550 ( .A(weight_1_bias_2[2]), .B(n36153), .Y(n36143) );
  OAI2BB1XL U37551 ( .A0N(weight_1_bias_3[2]), .A1N(n36155), .B0(n36143), .Y(
        n14098) );
  NAND2XL U37552 ( .A(weight_1_bias_1[2]), .B(n36153), .Y(n36144) );
  OAI2BB1XL U37553 ( .A0N(weight_1_bias_2[2]), .A1N(n36155), .B0(n36144), .Y(
        n14097) );
  OAI2BB2XL U37554 ( .B0(n36145), .B1(n36153), .A0N(weight_1_bias_3[3]), .A1N(
        n36153), .Y(n14096) );
  NAND2XL U37555 ( .A(weight_1_bias_2[3]), .B(n36153), .Y(n36146) );
  OAI2BB1XL U37556 ( .A0N(weight_1_bias_3[3]), .A1N(n36155), .B0(n36146), .Y(
        n14095) );
  NAND2XL U37557 ( .A(weight_1_bias_1[3]), .B(n36153), .Y(n36147) );
  OAI2BB1XL U37558 ( .A0N(weight_1_bias_2[3]), .A1N(n36155), .B0(n36147), .Y(
        n14094) );
  OAI2BB2XL U37559 ( .B0(n36148), .B1(n36153), .A0N(weight_1_bias_3[4]), .A1N(
        n36153), .Y(n14093) );
  NAND2XL U37560 ( .A(weight_1_bias_2[4]), .B(n36153), .Y(n36149) );
  OAI2BB1XL U37561 ( .A0N(weight_1_bias_3[4]), .A1N(n36155), .B0(n36149), .Y(
        n14092) );
  NAND2XL U37562 ( .A(weight_1_bias_1[4]), .B(n36153), .Y(n36150) );
  OAI2BB1XL U37563 ( .A0N(weight_1_bias_2[4]), .A1N(n36155), .B0(n36150), .Y(
        n14091) );
  OAI2BB2XL U37564 ( .B0(n36151), .B1(n36153), .A0N(weight_1_bias_3[5]), .A1N(
        n36153), .Y(n14090) );
  NAND2XL U37565 ( .A(weight_1_bias_2[5]), .B(n36153), .Y(n36152) );
  OAI2BB1XL U37566 ( .A0N(weight_1_bias_3[5]), .A1N(n36155), .B0(n36152), .Y(
        n14089) );
  NAND2XL U37567 ( .A(weight_1_bias_1[5]), .B(n36153), .Y(n36154) );
  OAI2BB1XL U37568 ( .A0N(weight_1_bias_2[5]), .A1N(n36155), .B0(n36154), .Y(
        n14088) );
  INVXL U37569 ( .A(affine_2[21]), .Y(n36219) );
  INVXL U37570 ( .A(affine_2[4]), .Y(n36177) );
  INVXL U37571 ( .A(affine_2[19]), .Y(n36160) );
  INVXL U37572 ( .A(affine_2[2]), .Y(n36174) );
  INVXL U37573 ( .A(affine_2[17]), .Y(n36156) );
  OAI2BB1XL U37574 ( .A0N(n36156), .A1N(affine_2[1]), .B0(affine_2[16]), .Y(
        n36157) );
  OAI22XL U37575 ( .A0(affine_2[0]), .A1(n36157), .B0(n36156), .B1(affine_2[1]), .Y(n36158) );
  AOI222XL U37576 ( .A0(affine_2[18]), .A1(n36174), .B0(affine_2[18]), .B1(
        n36158), .C0(n36174), .C1(n36158), .Y(n36159) );
  AOI222XL U37577 ( .A0(affine_2[3]), .A1(n36160), .B0(affine_2[3]), .B1(
        n36159), .C0(n36160), .C1(n36159), .Y(n36161) );
  AOI222XL U37578 ( .A0(affine_2[20]), .A1(n36177), .B0(affine_2[20]), .B1(
        n36161), .C0(n36177), .C1(n36161), .Y(n36162) );
  AOI222XL U37579 ( .A0(affine_2[5]), .A1(n36219), .B0(affine_2[5]), .B1(
        n36162), .C0(n36219), .C1(n36162), .Y(n36163) );
  INVXL U37580 ( .A(affine_2[6]), .Y(n36179) );
  AOI222XL U37581 ( .A0(affine_2[22]), .A1(n36163), .B0(affine_2[22]), .B1(
        n36179), .C0(n36163), .C1(n36179), .Y(n36164) );
  INVXL U37582 ( .A(affine_2[23]), .Y(n36224) );
  AOI222XL U37583 ( .A0(affine_2[7]), .A1(n36164), .B0(affine_2[7]), .B1(
        n36224), .C0(n36164), .C1(n36224), .Y(n36166) );
  INVXL U37584 ( .A(affine_2[8]), .Y(n36165) );
  AOI222XL U37585 ( .A0(affine_2[24]), .A1(n36166), .B0(affine_2[24]), .B1(
        n36165), .C0(n36166), .C1(n36165), .Y(n36167) );
  INVXL U37586 ( .A(affine_2[25]), .Y(n36225) );
  AOI222XL U37587 ( .A0(affine_2[9]), .A1(n36167), .B0(affine_2[9]), .B1(
        n36225), .C0(n36167), .C1(n36225), .Y(n36170) );
  AOI2BB1XL U37588 ( .A0N(affine_2[26]), .A1N(n36170), .B0(affine_2[10]), .Y(
        n36168) );
  AOI211XL U37589 ( .A0(n36170), .A1(affine_2[26]), .B0(n36169), .C0(n36168), 
        .Y(n36206) );
  INVXL U37590 ( .A(affine_2[12]), .Y(n36190) );
  INVXL U37591 ( .A(affine_2[15]), .Y(n36194) );
  AOI22XL U37592 ( .A0(affine_2[11]), .A1(DP_OP_5170J1_126_4278_n31), .B0(
        affine_2[31]), .B1(n36194), .Y(n36171) );
  INVXL U37593 ( .A(affine_2[30]), .Y(n36237) );
  AOI22XL U37594 ( .A0(affine_2[13]), .A1(n28394), .B0(affine_2[14]), .B1(
        n36237), .Y(n36196) );
  OAI211XL U37595 ( .A0(affine_2[28]), .A1(n36190), .B0(n36171), .C0(n36196), 
        .Y(n36205) );
  INVXL U37596 ( .A(affine_2[10]), .Y(n36188) );
  INVXL U37597 ( .A(affine_2[41]), .Y(n36208) );
  INVXL U37598 ( .A(affine_2[37]), .Y(n36215) );
  INVXL U37599 ( .A(affine_2[35]), .Y(n36213) );
  INVXL U37600 ( .A(affine_2[33]), .Y(n36209) );
  OAI2BB1XL U37601 ( .A0N(n36209), .A1N(affine_2[1]), .B0(affine_2[32]), .Y(
        n36172) );
  OAI22XL U37602 ( .A0(affine_2[0]), .A1(n36172), .B0(n36209), .B1(affine_2[1]), .Y(n36173) );
  AOI222XL U37603 ( .A0(affine_2[34]), .A1(n36174), .B0(affine_2[34]), .B1(
        n36173), .C0(n36174), .C1(n36173), .Y(n36175) );
  AOI222XL U37604 ( .A0(affine_2[3]), .A1(n36213), .B0(affine_2[3]), .B1(
        n36175), .C0(n36213), .C1(n36175), .Y(n36176) );
  AOI222XL U37605 ( .A0(affine_2[36]), .A1(n36177), .B0(affine_2[36]), .B1(
        n36176), .C0(n36177), .C1(n36176), .Y(n36178) );
  AOI222XL U37606 ( .A0(affine_2[5]), .A1(n36215), .B0(affine_2[5]), .B1(
        n36178), .C0(n36215), .C1(n36178), .Y(n36180) );
  AOI222XL U37607 ( .A0(affine_2[38]), .A1(n36180), .B0(affine_2[38]), .B1(
        n36179), .C0(n36180), .C1(n36179), .Y(n36182) );
  INVXL U37608 ( .A(affine_2[39]), .Y(n36181) );
  AOI222XL U37609 ( .A0(affine_2[7]), .A1(n36182), .B0(affine_2[7]), .B1(
        n36181), .C0(n36182), .C1(n36181), .Y(n36185) );
  NAND2XL U37610 ( .A(affine_2[9]), .B(n36208), .Y(n36184) );
  OAI2BB1XL U37611 ( .A0N(n36185), .A1N(affine_2[40]), .B0(affine_2[8]), .Y(
        n36183) );
  OAI211XL U37612 ( .A0(n36185), .A1(affine_2[40]), .B0(n36184), .C0(n36183), 
        .Y(n36186) );
  OAI21XL U37613 ( .A0(affine_2[9]), .A1(n36208), .B0(n36186), .Y(n36187) );
  AOI222XL U37614 ( .A0(affine_2[42]), .A1(n36188), .B0(affine_2[42]), .B1(
        n36187), .C0(n36188), .C1(n36187), .Y(n36189) );
  AOI222XL U37615 ( .A0(affine_2[11]), .A1(n36189), .B0(affine_2[11]), .B1(
        DP_OP_5169J1_125_4278_n31), .C0(n36189), .C1(DP_OP_5169J1_125_4278_n31), .Y(n36191) );
  AOI222XL U37616 ( .A0(affine_2[44]), .A1(n36191), .B0(affine_2[44]), .B1(
        n36190), .C0(n36191), .C1(n36190), .Y(n36193) );
  INVXL U37617 ( .A(affine_2[14]), .Y(n36195) );
  OAI2BB2XL U37618 ( .B0(affine_2[46]), .B1(n36195), .A0N(n28207), .A1N(
        affine_2[13]), .Y(n36192) );
  AOI221XL U37619 ( .A0(affine_2[13]), .A1(n36193), .B0(n28207), .B1(n36193), 
        .C0(n36192), .Y(n36203) );
  NAND2XL U37620 ( .A(affine_2[47]), .B(n36194), .Y(n36202) );
  OAI2BB2XL U37621 ( .B0(affine_2[47]), .B1(n36194), .A0N(n36195), .A1N(
        affine_2[46]), .Y(n36201) );
  INVXL U37622 ( .A(affine_2[31]), .Y(n36238) );
  INVXL U37623 ( .A(affine_2[28]), .Y(n36233) );
  OAI22XL U37624 ( .A0(affine_2[13]), .A1(n28394), .B0(affine_2[12]), .B1(
        n36233), .Y(n36197) );
  AOI222XL U37625 ( .A0(n36238), .A1(affine_2[15]), .B0(n36197), .B1(n36196), 
        .C0(n36195), .C1(affine_2[30]), .Y(n36198) );
  AOI221XL U37626 ( .A0(n36203), .A1(n36202), .B0(n36201), .B1(n36202), .C0(
        n36200), .Y(n36204) );
  OAI211XL U37627 ( .A0(n36206), .A1(n36205), .B0(n36207), .C0(n36204), .Y(
        n36242) );
  OAI2BB1XL U37628 ( .A0N(n36207), .A1N(number_2), .B0(n36242), .Y(n14087) );
  INVXL U37629 ( .A(affine_2[26]), .Y(n36231) );
  OAI2BB2XL U37630 ( .B0(affine_2[25]), .B1(n36208), .A0N(n36231), .A1N(
        affine_2[42]), .Y(n36230) );
  INVXL U37631 ( .A(affine_2[38]), .Y(n36222) );
  OAI2BB1XL U37632 ( .A0N(n36209), .A1N(affine_2[17]), .B0(affine_2[32]), .Y(
        n36210) );
  OAI22XL U37633 ( .A0(affine_2[16]), .A1(n36210), .B0(n36209), .B1(
        affine_2[17]), .Y(n36212) );
  INVXL U37634 ( .A(affine_2[18]), .Y(n36211) );
  AOI222XL U37635 ( .A0(affine_2[34]), .A1(n36212), .B0(affine_2[34]), .B1(
        n36211), .C0(n36212), .C1(n36211), .Y(n36214) );
  AOI222XL U37636 ( .A0(affine_2[19]), .A1(n36214), .B0(affine_2[19]), .B1(
        n36213), .C0(n36214), .C1(n36213), .Y(n36218) );
  AOI2BB1XL U37637 ( .A0N(affine_2[36]), .A1N(n36218), .B0(affine_2[20]), .Y(
        n36216) );
  AOI211XL U37638 ( .A0(n36218), .A1(affine_2[36]), .B0(n36217), .C0(n36216), 
        .Y(n36221) );
  OAI2BB2XL U37639 ( .B0(affine_2[37]), .B1(n36219), .A0N(n36222), .A1N(
        affine_2[22]), .Y(n36220) );
  OAI22XL U37640 ( .A0(affine_2[22]), .A1(n36222), .B0(n36221), .B1(n36220), 
        .Y(n36223) );
  AOI222XL U37641 ( .A0(affine_2[39]), .A1(n36224), .B0(affine_2[39]), .B1(
        n36223), .C0(n36224), .C1(n36223), .Y(n36228) );
  AOI2BB1XL U37642 ( .A0N(affine_2[24]), .A1N(n36228), .B0(affine_2[40]), .Y(
        n36226) );
  AOI211XL U37643 ( .A0(n36228), .A1(affine_2[24]), .B0(n36227), .C0(n36226), 
        .Y(n36229) );
  OAI22XL U37644 ( .A0(affine_2[42]), .A1(n36231), .B0(n36230), .B1(n36229), 
        .Y(n36232) );
  AOI222XL U37645 ( .A0(affine_2[27]), .A1(DP_OP_5169J1_125_4278_n31), .B0(
        affine_2[27]), .B1(n36232), .C0(DP_OP_5169J1_125_4278_n31), .C1(n36232), .Y(n36234) );
  AOI222XL U37646 ( .A0(affine_2[44]), .A1(n36234), .B0(affine_2[44]), .B1(
        n36233), .C0(n36234), .C1(n36233), .Y(n36235) );
  AOI222XL U37647 ( .A0(affine_2[29]), .A1(n28207), .B0(affine_2[29]), .B1(
        n36235), .C0(n28207), .C1(n36235), .Y(n36236) );
  AOI222XL U37648 ( .A0(affine_2[46]), .A1(n36237), .B0(affine_2[46]), .B1(
        n36236), .C0(n36237), .C1(n36236), .Y(n36239) );
  AOI222XL U37649 ( .A0(affine_2[47]), .A1(n36239), .B0(affine_2[47]), .B1(
        n36238), .C0(n36239), .C1(n36238), .Y(n36241) );
  AOI21XL U37650 ( .A0(n36242), .A1(n36241), .B0(number_6), .Y(n36240) );
  NOR2BXL U37651 ( .AN(n36242), .B(n36241), .Y(n36243) );
  AOI2BB1XL U37652 ( .A0N(n36243), .A1N(number_4), .B0(n36250), .Y(n14085) );
  CMPR42X1 U37653 ( .A(affine_2[20]), .B(DP_OP_5170J1_126_4278_n89), .C(
        DP_OP_5170J1_126_4278_n107), .D(DP_OP_5170J1_126_4278_n98), .ICI(
        DP_OP_5170J1_126_4278_n67), .S(DP_OP_5170J1_126_4278_n64), .ICO(
        DP_OP_5170J1_126_4278_n62), .CO(DP_OP_5170J1_126_4278_n63) );
endmodule

